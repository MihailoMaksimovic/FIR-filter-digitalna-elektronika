magic
tech sky130A
timestamp 1693223098
<< nwell >>
rect -120 -25 295 115
<< nmos >>
rect 0 -300 15 -200
rect 65 -300 80 -200
rect 210 -300 225 -200
<< pmos >>
rect 0 -5 15 95
rect 65 -5 80 95
rect 210 -5 225 95
<< ndiff >>
rect -50 -215 0 -200
rect -50 -285 -35 -215
rect -15 -285 0 -215
rect -50 -300 0 -285
rect 15 -215 65 -200
rect 15 -285 30 -215
rect 50 -285 65 -215
rect 15 -300 65 -285
rect 80 -215 130 -200
rect 80 -285 95 -215
rect 115 -285 130 -215
rect 80 -300 130 -285
rect 160 -215 210 -200
rect 160 -285 175 -215
rect 195 -285 210 -215
rect 160 -300 210 -285
rect 225 -215 275 -200
rect 225 -285 240 -215
rect 260 -285 275 -215
rect 225 -300 275 -285
<< pdiff >>
rect -50 80 0 95
rect -50 10 -35 80
rect -15 10 0 80
rect -50 -5 0 10
rect 15 80 65 95
rect 15 10 30 80
rect 50 10 65 80
rect 15 -5 65 10
rect 80 80 130 95
rect 80 10 95 80
rect 115 10 130 80
rect 80 -5 130 10
rect 160 80 210 95
rect 160 10 175 80
rect 195 10 210 80
rect 160 -5 210 10
rect 225 80 275 95
rect 225 10 240 80
rect 260 10 275 80
rect 225 -5 275 10
<< ndiffc >>
rect -35 -285 -15 -215
rect 30 -285 50 -215
rect 95 -285 115 -215
rect 175 -285 195 -215
rect 240 -285 260 -215
<< pdiffc >>
rect -35 10 -15 80
rect 30 10 50 80
rect 95 10 115 80
rect 175 10 195 80
rect 240 10 260 80
<< psubdiff >>
rect -100 -215 -50 -200
rect -100 -285 -85 -215
rect -65 -285 -50 -215
rect -100 -300 -50 -285
<< nsubdiff >>
rect -100 80 -50 95
rect -100 10 -85 80
rect -65 10 -50 80
rect -100 -5 -50 10
<< psubdiffcont >>
rect -85 -285 -65 -215
<< nsubdiffcont >>
rect -85 10 -65 80
<< poly >>
rect 0 95 15 110
rect 65 95 80 110
rect 210 95 225 110
rect 0 -25 15 -5
rect -25 -35 15 -25
rect -25 -55 -15 -35
rect 5 -55 15 -35
rect -25 -65 15 -55
rect 0 -200 15 -65
rect 65 -100 80 -5
rect 210 -25 225 -5
rect 185 -35 225 -25
rect 185 -55 195 -35
rect 215 -55 225 -35
rect 185 -65 225 -55
rect 40 -110 80 -100
rect 40 -130 50 -110
rect 70 -130 80 -110
rect 40 -140 80 -130
rect 65 -200 80 -140
rect 210 -200 225 -65
rect 0 -315 15 -300
rect 65 -315 80 -300
rect 210 -315 225 -300
<< polycont >>
rect -15 -55 5 -35
rect 195 -55 215 -35
rect 50 -130 70 -110
<< locali >>
rect -95 80 -5 90
rect -95 10 -85 80
rect -65 10 -35 80
rect -15 10 -5 80
rect -95 0 -5 10
rect 20 80 60 90
rect 20 10 30 80
rect 50 10 60 80
rect 20 0 60 10
rect 85 80 125 90
rect 85 10 95 80
rect 115 10 125 80
rect 85 0 125 10
rect 160 80 205 90
rect 160 10 175 80
rect 195 10 205 80
rect 160 0 205 10
rect 230 80 270 90
rect 230 10 240 80
rect 260 10 270 80
rect 230 0 270 10
rect 40 -25 60 0
rect 250 -25 270 0
rect -120 -35 15 -25
rect -120 -45 -15 -35
rect -25 -55 -15 -45
rect 5 -55 15 -35
rect 40 -35 225 -25
rect 40 -45 195 -35
rect -25 -65 15 -55
rect -120 -110 80 -100
rect -120 -120 50 -110
rect 40 -130 50 -120
rect 70 -130 80 -110
rect 40 -140 80 -130
rect 105 -205 125 -45
rect 185 -55 195 -45
rect 215 -55 225 -35
rect 185 -65 225 -55
rect 250 -45 295 -25
rect 250 -205 270 -45
rect -95 -215 -5 -205
rect -95 -285 -85 -215
rect -65 -285 -35 -215
rect -15 -285 -5 -215
rect -95 -295 -5 -285
rect 20 -215 60 -205
rect 20 -285 30 -215
rect 50 -285 60 -215
rect 20 -295 60 -285
rect 85 -215 125 -205
rect 85 -285 95 -215
rect 115 -285 125 -215
rect 85 -295 125 -285
rect 160 -215 205 -205
rect 160 -285 175 -215
rect 195 -285 205 -215
rect 160 -295 205 -285
rect 230 -215 270 -205
rect 230 -285 240 -215
rect 260 -285 270 -215
rect 230 -295 270 -285
<< viali >>
rect -85 10 -65 80
rect -35 10 -15 80
rect 95 10 115 80
rect 175 10 195 80
rect -85 -285 -65 -215
rect -35 -285 -15 -215
rect 175 -285 195 -215
<< metal1 >>
rect -120 80 295 95
rect -120 10 -85 80
rect -65 10 -35 80
rect -15 10 95 80
rect 115 10 175 80
rect 195 10 295 80
rect -120 -5 295 10
rect -120 -215 295 -200
rect -120 -285 -85 -215
rect -65 -285 -35 -215
rect -15 -285 175 -215
rect 195 -285 295 -215
rect -120 -300 295 -285
<< labels >>
rlabel locali -120 -35 -120 -35 7 A
port 1 w
rlabel locali -120 -110 -120 -110 7 B
port 2 w
rlabel metal1 -120 -250 -120 -250 7 VN
port 5 w
rlabel metal1 -120 45 -120 45 7 VP
port 4 w
rlabel locali 295 -35 295 -35 3 X
port 3 e
<< end >>
