** sch_path: /home/mihailo/projekat_sky130/projekat_layout/fa_8bits/FA_8bits.sch
**.subckt FA_8bits A0 B0 A1 B1 S0 S1 VP VN Cin_first A2 B2 S2 A3 B3 S3 A4 B4 S4 A5 B5 S5 A6 B6 S6 S7
*+ A7 B7 S8
*.ipin A0
*.ipin B0
*.ipin A1
*.ipin B1
*.opin S0
*.opin S1
*.iopin VP
*.iopin VN
*.ipin Cin_first
*.ipin A2
*.ipin B2
*.opin S2
*.ipin A3
*.ipin B3
*.opin S3
*.ipin A4
*.ipin B4
*.opin S4
*.ipin A5
*.ipin B5
*.opin S5
*.ipin A6
*.ipin B6
*.opin S6
*.opin S7
*.ipin A7
*.ipin B7
*.opin S8
X1 A0 B0 Cin_first net1 S0 VP VN FA
X2 A1 B1 net1 net2 S1 VP VN FA
X3 A2 B2 net2 net3 S2 VP VN FA
X4 A3 B3 net3 net4 S3 VP VN FA
X5 A4 B4 net4 net5 S4 VP VN FA
X6 A5 B5 net5 net6 S5 VP VN FA
X7 A6 B6 net6 net7 S6 VP VN FA
X8 A7 B7 net7 S8 S7 VP VN FA
**.ends

* expanding   symbol:  /home/mihailo/projekat_sky130/projekat_layout/fa/FA.sym # of pins=7
** sym_path: /home/mihailo/projekat_sky130/projekat_layout/fa/FA.sym
** sch_path: /home/mihailo/projekat_sky130/projekat_layout/fa/FA.sch
.subckt FA A B Cin Out Sum VP VN
*.ipin A
*.opin Sum
*.iopin VP
*.iopin VN
*.opin Out
*.ipin B
*.ipin Cin
X4 A B VN VP net1 XOR
X5 Cin net1 VN VP Sum XOR
X1 Cin net1 net3 VP VN AND
X2 A B net2 VP VN AND
X3 net3 net2 Out VP VN OR
.ends


* expanding   symbol:  /home/mihailo/projekat_sky130/projekat_layout/xor/XOR.sym # of pins=5
** sym_path: /home/mihailo/projekat_sky130/projekat_layout/xor/XOR.sym
** sch_path: /home/mihailo/projekat_sky130/projekat_layout/xor/XOR.sch
.subckt XOR A B VN VP X
*.ipin A
*.ipin B
*.opin X
*.iopin VN
*.iopin VP
X1 B net3 net1 VP VN AND
X2 net4 A net2 VP VN AND
X3 net1 net2 X VP VN OR
X4 A net3 VP VN invertor
X5 B net4 VP VN invertor
.ends


* expanding   symbol:  /home/mihailo/projekat_sky130/projekat_layout/and/AND.sym # of pins=5
** sym_path: /home/mihailo/projekat_sky130/projekat_layout/and/AND.sym
** sch_path: /home/mihailo/projekat_sky130/projekat_layout/and/AND.sch
.subckt AND A B X VP VN
*.ipin A
*.ipin B
*.iopin VN
*.iopin VP
*.opin X
XM1 net1 A net2 VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 B VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 B VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 X net1 VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 X net1 VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /home/mihailo/projekat_sky130/projekat_layout/or/OR.sym # of pins=5
** sym_path: /home/mihailo/projekat_sky130/projekat_layout/or/OR.sym
** sch_path: /home/mihailo/projekat_sky130/projekat_layout/or/OR.sch
.subckt OR A B X VP VN
*.opin X
*.ipin A
*.ipin B
*.iopin VP
*.iopin VN
XM1 net2 A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 B net1 VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 B VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 X net2 VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 X net2 VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /home/mihailo/projekat_sky130/projekat_layout/invertor/invertor.sym # of
*+ pins=4
** sym_path: /home/mihailo/projekat_sky130/projekat_layout/invertor/invertor.sym
** sch_path: /home/mihailo/projekat_sky130/projekat_layout/invertor/invertor.sch
.subckt invertor A Y VP VN
*.iopin VP
*.iopin VN
*.ipin A
*.opin Y
XM1 Y A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
