magic
tech sky130A
timestamp 1693914941
<< nwell >>
rect 2420 1220 2605 1360
rect 4915 1215 5090 1355
rect 7410 1210 7570 1350
rect 9900 1210 10060 1350
rect 12380 1210 12560 1350
rect 14880 1210 15040 1350
rect 17370 1210 17530 1350
<< poly >>
rect 2405 1725 2445 1735
rect 2405 1705 2415 1725
rect 2435 1705 2445 1725
rect 2405 1695 2445 1705
rect 2430 850 2445 1695
rect 4895 1720 4935 1730
rect 4895 1700 4905 1720
rect 4925 1700 4935 1720
rect 4895 1690 4935 1700
rect 7385 1720 7425 1730
rect 7385 1700 7395 1720
rect 7415 1700 7425 1720
rect 7385 1690 7425 1700
rect 9875 1720 9915 1730
rect 9875 1700 9885 1720
rect 9905 1700 9915 1720
rect 9875 1690 9915 1700
rect 12370 1720 12410 1730
rect 12370 1700 12380 1720
rect 12400 1700 12410 1720
rect 12370 1690 12410 1700
rect 14855 1715 14895 1725
rect 14855 1695 14865 1715
rect 14885 1695 14895 1715
rect 2405 840 2445 850
rect 4920 845 4935 1690
rect 2405 820 2415 840
rect 2435 820 2445 840
rect 2405 810 2445 820
rect 4895 835 4935 845
rect 7410 840 7425 1690
rect 9900 840 9915 1690
rect 4895 815 4905 835
rect 4925 815 4935 835
rect 4895 805 4935 815
rect 7385 830 7425 840
rect 7385 810 7395 830
rect 7415 810 7425 830
rect 7385 800 7425 810
rect 9875 830 9915 840
rect 12390 835 12405 1690
rect 14855 1685 14895 1695
rect 17345 1720 17385 1730
rect 17345 1700 17355 1720
rect 17375 1700 17385 1720
rect 17345 1690 17385 1700
rect 14880 840 14895 1685
rect 17370 840 17385 1690
rect 9875 810 9885 830
rect 9905 810 9915 830
rect 9875 800 9915 810
rect 12365 825 12405 835
rect 12365 805 12375 825
rect 12395 805 12405 825
rect 12365 795 12405 805
rect 14855 830 14895 840
rect 14855 810 14865 830
rect 14885 810 14895 830
rect 14855 800 14895 810
rect 17350 830 17390 840
rect 17350 810 17360 830
rect 17380 810 17390 830
rect 17350 800 17390 810
<< polycont >>
rect 2415 1705 2435 1725
rect 4905 1700 4925 1720
rect 7395 1700 7415 1720
rect 9885 1700 9905 1720
rect 12380 1700 12400 1720
rect 14865 1695 14885 1715
rect 2415 820 2435 840
rect 4905 815 4925 835
rect 7395 810 7415 830
rect 17355 1700 17375 1720
rect 9885 810 9905 830
rect 12375 805 12395 825
rect 14865 810 14885 830
rect 17360 810 17380 830
<< locali >>
rect 2405 1725 2565 1735
rect 2405 1705 2415 1725
rect 2435 1715 2565 1725
rect 4895 1720 5055 1730
rect 2435 1705 2445 1715
rect 2405 1695 2445 1705
rect 4895 1700 4905 1720
rect 4925 1710 5055 1720
rect 7385 1720 7545 1730
rect 4925 1700 4935 1710
rect 4895 1690 4935 1700
rect 5055 1690 5060 1710
rect 7385 1700 7395 1720
rect 7415 1710 7545 1720
rect 9875 1720 10035 1730
rect 7415 1700 7425 1710
rect 7385 1690 7425 1700
rect 9875 1700 9885 1720
rect 9905 1710 10035 1720
rect 12370 1720 12530 1730
rect 9905 1700 9920 1710
rect 9875 1690 9920 1700
rect 12370 1700 12380 1720
rect 12400 1710 12530 1720
rect 14855 1715 15015 1730
rect 12400 1700 12415 1710
rect 12370 1690 12415 1700
rect 14855 1695 14865 1715
rect 14885 1710 15015 1715
rect 17345 1720 17505 1730
rect 14885 1695 14895 1710
rect 14855 1685 14895 1695
rect 17345 1700 17355 1720
rect 17375 1710 17505 1720
rect 17375 1700 17385 1710
rect 17345 1690 17385 1700
rect 4915 1195 4935 1215
rect 2405 840 2445 850
rect 2405 830 2415 840
rect 980 820 2415 830
rect 2435 820 2445 840
rect 4895 835 4935 845
rect 4895 825 4905 835
rect 980 810 2445 820
rect 3470 815 4905 825
rect 4925 815 4935 835
rect 7385 830 7425 840
rect 7385 820 7395 830
rect 980 615 1000 810
rect 3470 805 4935 815
rect 5960 810 7395 820
rect 7415 810 7425 830
rect 9875 830 9915 840
rect 9875 820 9885 830
rect 3470 630 3490 805
rect 3445 610 3490 630
rect 5960 800 7425 810
rect 8450 810 9885 820
rect 9905 810 9915 830
rect 12365 825 12405 835
rect 12365 815 12375 825
rect 8450 800 9915 810
rect 10940 805 12375 815
rect 12395 805 12405 825
rect 14855 830 14895 840
rect 14855 820 14865 830
rect 5960 605 5980 800
rect 8450 605 8470 800
rect 10940 795 12405 805
rect 13430 810 14865 820
rect 14885 810 14895 830
rect 17350 830 17390 840
rect 17350 820 17360 830
rect 13430 800 14895 810
rect 15920 810 17360 820
rect 17380 810 17390 830
rect 15920 800 17390 810
rect 10940 605 10960 795
rect 13430 605 13450 800
rect 15920 605 15945 800
<< metal1 >>
rect 2420 945 2665 1045
rect 4910 940 5155 1040
rect 7405 935 7635 1035
rect 9890 935 10140 1035
rect 12385 935 12625 1035
rect 14875 935 15115 1035
rect 17365 935 17600 1035
use fa  fa_0
timestamp 1693913107
transform 1 0 90 0 1 930
box -140 -930 2340 975
use fa  fa_1
timestamp 1693913107
transform 1 0 2580 0 1 925
box -140 -930 2340 975
use fa  fa_2
timestamp 1693913107
transform 1 0 5070 0 1 920
box -140 -930 2340 975
use fa  fa_3
timestamp 1693913107
transform 1 0 7560 0 1 920
box -140 -930 2340 975
use fa  fa_4
timestamp 1693913107
transform 1 0 10050 0 1 920
box -140 -930 2340 975
use fa  fa_5
timestamp 1693913107
transform 1 0 12540 0 1 920
box -140 -930 2340 975
use fa  fa_6
timestamp 1693913107
transform 1 0 15030 0 1 920
box -140 -930 2340 975
use fa  fa_7
timestamp 1693913107
transform 1 0 17520 0 1 920
box -140 -930 2340 975
<< end >>
