magic
tech sky130A
timestamp 1693949129
<< nwell >>
rect 27860 1780 28190 1795
rect 27845 1675 28190 1780
rect 27860 1655 28190 1675
rect 27870 780 28180 885
rect 27870 -1705 28005 780
rect 27870 -1830 28190 -1705
rect 27945 -1845 28190 -1830
rect 27860 -5350 28190 -5335
rect 27845 -5455 28190 -5350
rect 27860 -5475 28190 -5455
rect 27910 -9365 28190 -9225
rect 27910 -12475 28025 -9365
rect 27860 -12490 28190 -12475
rect 27845 -12595 28190 -12490
rect 27860 -12615 28190 -12595
<< ndiff >>
rect 30365 -2155 30405 -2145
rect 30365 -2175 30375 -2155
rect 30395 -2175 30405 -2155
rect 30365 -2185 30405 -2175
rect 32855 -2155 32895 -2145
rect 32855 -2175 32865 -2155
rect 32885 -2175 32895 -2155
rect 32855 -2185 32895 -2175
rect 35345 -2155 35385 -2145
rect 35345 -2175 35355 -2155
rect 35375 -2175 35385 -2155
rect 35345 -2185 35385 -2175
rect 37835 -2155 37875 -2145
rect 37835 -2175 37845 -2155
rect 37865 -2175 37875 -2155
rect 37835 -2185 37875 -2175
rect 40325 -2155 40365 -2145
rect 40325 -2175 40335 -2155
rect 40355 -2175 40365 -2155
rect 40325 -2185 40365 -2175
rect 42815 -2155 42855 -2145
rect 42815 -2175 42825 -2155
rect 42845 -2175 42855 -2155
rect 42815 -2185 42855 -2175
rect 45305 -2155 45345 -2145
rect 45305 -2175 45315 -2155
rect 45335 -2175 45345 -2155
rect 45305 -2185 45345 -2175
rect 47795 -2155 47835 -2145
rect 47795 -2175 47805 -2155
rect 47825 -2175 47835 -2155
rect 47795 -2185 47835 -2175
rect 30365 -8155 30405 -8145
rect 30365 -8175 30375 -8155
rect 30395 -8175 30405 -8155
rect 30365 -8185 30405 -8175
rect 32855 -8155 32895 -8145
rect 32855 -8175 32865 -8155
rect 32885 -8175 32895 -8155
rect 32855 -8185 32895 -8175
rect 35345 -8155 35385 -8145
rect 35345 -8175 35355 -8155
rect 35375 -8175 35385 -8155
rect 35345 -8185 35385 -8175
rect 37835 -8155 37875 -8145
rect 37835 -8175 37845 -8155
rect 37865 -8175 37875 -8155
rect 37835 -8185 37875 -8175
rect 40325 -8155 40365 -8145
rect 40325 -8175 40335 -8155
rect 40355 -8175 40365 -8155
rect 40325 -8185 40365 -8175
rect 42815 -8155 42855 -8145
rect 42815 -8175 42825 -8155
rect 42845 -8175 42855 -8155
rect 42815 -8185 42855 -8175
rect 45305 -8155 45345 -8145
rect 45305 -8175 45315 -8155
rect 45335 -8175 45345 -8155
rect 45305 -8185 45345 -8175
rect 47795 -8155 47835 -8145
rect 47795 -8175 47805 -8155
rect 47825 -8175 47835 -8155
rect 47795 -8185 47835 -8175
<< ndiffc >>
rect 30375 -2175 30395 -2155
rect 32865 -2175 32885 -2155
rect 35355 -2175 35375 -2155
rect 37845 -2175 37865 -2155
rect 40335 -2175 40355 -2155
rect 42825 -2175 42845 -2155
rect 45315 -2175 45335 -2155
rect 47805 -2175 47825 -2155
rect 30375 -8175 30395 -8155
rect 32865 -8175 32885 -8155
rect 35355 -8175 35375 -8155
rect 37845 -8175 37865 -8155
rect 40335 -8175 40355 -8155
rect 42825 -8175 42845 -8155
rect 45315 -8175 45335 -8155
rect 47805 -8175 47825 -8155
<< poly >>
rect 125 6790 165 6800
rect 125 6770 135 6790
rect 155 6770 165 6790
rect 125 6760 165 6770
rect 1805 6790 1845 6800
rect 1805 6770 1815 6790
rect 1835 6770 1845 6790
rect 1805 6760 1845 6770
rect 2935 6790 2975 6800
rect 2935 6770 2945 6790
rect 2965 6770 2975 6790
rect 2935 6760 2975 6770
rect 4065 6790 4105 6800
rect 4065 6770 4075 6790
rect 4095 6770 4105 6790
rect 4065 6760 4105 6770
rect 5695 6790 5735 6800
rect 5695 6770 5705 6790
rect 5725 6770 5735 6790
rect 5695 6760 5735 6770
rect 6825 6790 6865 6800
rect 6825 6770 6835 6790
rect 6855 6770 6865 6790
rect 6825 6760 6865 6770
rect 125 6090 140 6760
rect 1125 6495 1165 6505
rect 1125 6475 1135 6495
rect 1155 6475 1165 6495
rect 1125 6465 1165 6475
rect 60 -550 75 1020
rect 125 -330 140 650
rect 1150 65 1165 6465
rect 1805 6090 1820 6760
rect 2935 6090 2950 6760
rect 4065 6090 4080 6760
rect 5060 6495 5100 6505
rect 5060 6475 5070 6495
rect 5090 6475 5100 6495
rect 5060 6465 5100 6475
rect 1125 55 1165 65
rect 1125 35 1135 55
rect 1155 35 1165 55
rect 1125 25 1165 35
rect 1190 5845 1230 5855
rect 1190 5825 1200 5845
rect 1220 5825 1230 5845
rect 1190 5815 1230 5825
rect 1190 0 1205 5815
rect 1250 4945 1290 4955
rect 1250 4925 1260 4945
rect 1280 4925 1290 4945
rect 1250 4915 1290 4925
rect 1165 -10 1205 0
rect 1165 -30 1175 -10
rect 1195 -30 1205 -10
rect 1165 -40 1205 -30
rect 1275 -60 1290 4915
rect 1320 4045 1360 4055
rect 1320 4025 1330 4045
rect 1350 4025 1360 4045
rect 1320 4015 1360 4025
rect 1275 -70 1315 -60
rect 1275 -90 1285 -70
rect 1305 -90 1315 -70
rect 1275 -100 1315 -90
rect 1345 -105 1360 4015
rect 1385 3145 1425 3155
rect 1385 3125 1395 3145
rect 1415 3125 1425 3145
rect 1385 3115 1425 3125
rect 1345 -115 1385 -105
rect 1345 -135 1355 -115
rect 1375 -135 1385 -115
rect 1345 -145 1385 -135
rect 1410 -150 1425 3115
rect 1450 2245 1490 2255
rect 1450 2225 1460 2245
rect 1480 2225 1490 2245
rect 1450 2215 1490 2225
rect 1410 -160 1450 -150
rect 1410 -180 1420 -160
rect 1440 -180 1450 -160
rect 1410 -190 1450 -180
rect 1475 -195 1490 2215
rect 1520 1345 1560 1355
rect 1520 1325 1530 1345
rect 1550 1325 1560 1345
rect 1520 1315 1560 1325
rect 1475 -205 1515 -195
rect 1475 -225 1485 -205
rect 1505 -225 1515 -205
rect 1475 -235 1515 -225
rect 1545 -240 1560 1315
rect 1615 605 1655 615
rect 1615 585 1625 605
rect 1645 585 1655 605
rect 1615 575 1655 585
rect 1545 -250 1585 -240
rect 1545 -270 1555 -250
rect 1575 -270 1585 -250
rect 1545 -280 1585 -270
rect 1615 -290 1630 575
rect 5085 455 5100 6465
rect 5695 6090 5710 6760
rect 6825 6080 6840 6760
rect 7845 6005 7885 6015
rect 7845 5985 7855 6005
rect 7875 5990 7885 6005
rect 7875 5985 8010 5990
rect 7845 5975 8010 5985
rect 5060 445 5100 455
rect 5060 425 5070 445
rect 5090 425 5100 445
rect 5060 415 5100 425
rect 5125 5845 5165 5855
rect 5125 5825 5135 5845
rect 5155 5825 5165 5845
rect 5125 5815 5165 5825
rect 5125 390 5140 5815
rect 5185 4945 5225 4955
rect 5185 4925 5195 4945
rect 5215 4925 5225 4945
rect 5185 4915 5225 4925
rect 5100 380 5140 390
rect 5100 360 5110 380
rect 5130 360 5140 380
rect 5100 350 5140 360
rect 5210 330 5225 4915
rect 5255 4045 5295 4055
rect 5255 4025 5265 4045
rect 5285 4025 5295 4045
rect 5255 4015 5295 4025
rect 5210 320 5250 330
rect 5210 300 5220 320
rect 5240 300 5250 320
rect 5210 290 5250 300
rect 5280 285 5295 4015
rect 5320 3145 5360 3155
rect 5320 3125 5330 3145
rect 5350 3125 5360 3145
rect 5320 3115 5360 3125
rect 5280 275 5320 285
rect 5280 255 5290 275
rect 5310 255 5320 275
rect 5280 245 5320 255
rect 5345 240 5360 3115
rect 5385 2245 5425 2255
rect 5385 2225 5395 2245
rect 5415 2225 5425 2245
rect 5385 2215 5425 2225
rect 5345 230 5385 240
rect 5345 210 5355 230
rect 5375 210 5385 230
rect 5345 200 5385 210
rect 5410 195 5425 2215
rect 7995 2145 8010 5975
rect 8040 5845 8080 5855
rect 8040 5825 8050 5845
rect 8070 5825 8080 5845
rect 8040 5815 8080 5825
rect 8040 2370 8055 5815
rect 8085 4945 8125 4955
rect 8085 4925 8095 4945
rect 8115 4925 8125 4945
rect 8085 4915 8125 4925
rect 8085 2410 8100 4915
rect 8135 4045 8175 4055
rect 8135 4025 8145 4045
rect 8165 4025 8175 4045
rect 8135 4015 8175 4025
rect 8135 2450 8150 4015
rect 8185 3145 8225 3155
rect 8185 3125 8195 3145
rect 8215 3125 8225 3145
rect 8185 3115 8225 3125
rect 8185 2490 8200 3115
rect 25915 3110 25955 3120
rect 25915 3090 25925 3110
rect 25945 3090 25955 3110
rect 25915 3080 25955 3090
rect 8375 2625 8415 2635
rect 8375 2605 8385 2625
rect 8405 2610 8415 2625
rect 8405 2605 25440 2610
rect 8375 2595 25440 2605
rect 8310 2585 8350 2595
rect 8310 2565 8320 2585
rect 8340 2570 8350 2585
rect 8340 2565 22950 2570
rect 8310 2555 22950 2565
rect 8245 2545 8285 2555
rect 8245 2525 8255 2545
rect 8275 2530 8285 2545
rect 8275 2525 20460 2530
rect 8245 2515 20460 2525
rect 8185 2475 17970 2490
rect 8135 2435 15480 2450
rect 8085 2395 12990 2410
rect 8040 2355 10500 2370
rect 10485 2140 10500 2355
rect 12975 2135 12990 2395
rect 15465 2135 15480 2435
rect 17955 2135 17970 2475
rect 20445 2135 20460 2515
rect 22935 2135 22950 2555
rect 25425 2135 25440 2595
rect 25915 2325 25930 3080
rect 25980 3060 26020 3070
rect 25980 3040 25990 3060
rect 26010 3040 26020 3060
rect 25980 3030 26020 3040
rect 25980 2370 25995 3030
rect 26050 3015 26090 3025
rect 26050 2995 26060 3015
rect 26080 2995 26090 3015
rect 26050 2985 26090 2995
rect 26050 2410 26065 2985
rect 26130 2965 26170 2975
rect 26130 2945 26140 2965
rect 26160 2945 26170 2965
rect 26130 2935 26170 2945
rect 26130 2450 26145 2935
rect 26195 2915 26235 2925
rect 26195 2895 26205 2915
rect 26225 2895 26235 2915
rect 26195 2885 26235 2895
rect 26195 2490 26210 2885
rect 26265 2870 26305 2880
rect 26265 2850 26275 2870
rect 26295 2850 26305 2870
rect 26265 2840 26305 2850
rect 26265 2530 26280 2840
rect 26335 2825 26375 2835
rect 26335 2805 26345 2825
rect 26365 2805 26375 2825
rect 26335 2795 26375 2805
rect 26335 2570 26350 2795
rect 27860 2625 27900 2635
rect 27860 2605 27870 2625
rect 27890 2610 27900 2625
rect 27890 2605 45515 2610
rect 27860 2595 45515 2605
rect 26335 2555 43025 2570
rect 26265 2515 40535 2530
rect 26195 2475 38045 2490
rect 26130 2435 35555 2450
rect 26050 2395 33065 2410
rect 25980 2355 30575 2370
rect 25915 2310 28085 2325
rect 28070 2150 28085 2310
rect 30560 2145 30575 2355
rect 33050 2140 33065 2395
rect 35540 2140 35555 2435
rect 38030 2140 38045 2475
rect 40520 2140 40535 2515
rect 43010 2140 43025 2555
rect 45500 2140 45515 2595
rect 5455 1345 5495 1355
rect 5455 1325 5465 1345
rect 5485 1325 5495 1345
rect 5455 1315 5495 1325
rect 30400 1345 30440 1355
rect 30400 1325 30410 1345
rect 30430 1325 30440 1345
rect 30400 1315 30440 1325
rect 5410 185 5450 195
rect 5410 165 5420 185
rect 5440 165 5450 185
rect 5410 155 5450 165
rect 5480 150 5495 1315
rect 5550 585 5590 595
rect 5550 565 5560 585
rect 5580 565 5590 585
rect 5550 555 5590 565
rect 5480 140 5520 150
rect 5480 120 5490 140
rect 5510 120 5520 140
rect 5480 110 5520 120
rect 5550 105 5565 555
rect 8010 435 8025 740
rect 10500 435 10515 735
rect 12990 435 13005 730
rect 15480 435 15495 730
rect 17970 435 17985 730
rect 20460 435 20475 730
rect 22950 435 22965 730
rect 25440 435 25455 730
rect 7985 425 8025 435
rect 7985 405 7995 425
rect 8015 405 8025 425
rect 7985 395 8025 405
rect 10475 425 10515 435
rect 10475 405 10485 425
rect 10505 405 10515 425
rect 10475 395 10515 405
rect 12965 425 13005 435
rect 12965 405 12975 425
rect 12995 405 13005 425
rect 12965 395 13005 405
rect 15455 425 15495 435
rect 15455 405 15465 425
rect 15485 405 15495 425
rect 15455 395 15495 405
rect 17945 425 17985 435
rect 17945 405 17955 425
rect 17975 405 17985 425
rect 17945 395 17985 405
rect 20435 425 20475 435
rect 20435 405 20445 425
rect 20465 405 20475 425
rect 20435 395 20475 405
rect 22925 425 22965 435
rect 22925 405 22935 425
rect 22955 405 22965 425
rect 22925 395 22965 405
rect 25415 425 25455 435
rect 25415 405 25425 425
rect 25445 405 25455 425
rect 25415 395 25455 405
rect 28085 390 28100 745
rect 28060 380 28100 390
rect 28060 360 28070 380
rect 28090 360 28100 380
rect 28060 350 28100 360
rect 5550 95 5590 105
rect 5550 75 5560 95
rect 5580 75 5590 95
rect 5550 65 5590 75
rect 1615 -300 1655 -290
rect 1615 -320 1625 -300
rect 1645 -320 1655 -300
rect 1615 -330 1655 -320
rect 125 -340 165 -330
rect 125 -360 135 -340
rect 155 -360 165 -340
rect 125 -370 165 -360
rect 1255 -340 1295 -330
rect 1255 -360 1265 -340
rect 1285 -360 1295 -340
rect 1255 -370 1295 -360
rect 2935 -340 2975 -330
rect 2935 -360 2945 -340
rect 2965 -360 2975 -340
rect 2935 -370 2975 -360
rect 4065 -340 4105 -330
rect 4065 -360 4075 -340
rect 4095 -360 4105 -340
rect 4065 -370 4105 -360
rect 5170 -340 5210 -330
rect 5170 -360 5180 -340
rect 5200 -360 5210 -340
rect 5170 -370 5210 -360
rect 125 -1040 140 -370
rect 1255 -1040 1270 -370
rect 2250 -635 2290 -625
rect 2250 -655 2260 -635
rect 2280 -655 2290 -635
rect 2250 -665 2290 -655
rect 60 -7690 75 -6105
rect 125 -7470 140 -6480
rect 2275 -7065 2290 -665
rect 2935 -1040 2950 -370
rect 4065 -1040 4080 -370
rect 5195 -1040 5210 -370
rect 6825 -340 6865 -330
rect 6825 -360 6835 -340
rect 6855 -360 6865 -340
rect 6825 -370 6865 -360
rect 6185 -635 6225 -625
rect 6185 -655 6195 -635
rect 6215 -655 6225 -635
rect 6185 -665 6225 -655
rect 2250 -7075 2290 -7065
rect 2250 -7095 2260 -7075
rect 2280 -7095 2290 -7075
rect 2250 -7105 2290 -7095
rect 2315 -1285 2355 -1275
rect 2315 -1305 2325 -1285
rect 2345 -1305 2355 -1285
rect 2315 -1315 2355 -1305
rect 2315 -7130 2330 -1315
rect 2375 -2185 2415 -2175
rect 2375 -2205 2385 -2185
rect 2405 -2205 2415 -2185
rect 2375 -2215 2415 -2205
rect 2290 -7140 2330 -7130
rect 2290 -7160 2300 -7140
rect 2320 -7160 2330 -7140
rect 2290 -7170 2330 -7160
rect 2400 -7190 2415 -2215
rect 2445 -3085 2485 -3075
rect 2445 -3105 2455 -3085
rect 2475 -3105 2485 -3085
rect 2445 -3115 2485 -3105
rect 2400 -7200 2440 -7190
rect 2400 -7220 2410 -7200
rect 2430 -7220 2440 -7200
rect 2400 -7230 2440 -7220
rect 2470 -7235 2485 -3115
rect 2510 -3985 2550 -3975
rect 2510 -4005 2520 -3985
rect 2540 -4005 2550 -3985
rect 2510 -4015 2550 -4005
rect 2470 -7245 2510 -7235
rect 2470 -7265 2480 -7245
rect 2500 -7265 2510 -7245
rect 2470 -7275 2510 -7265
rect 2535 -7280 2550 -4015
rect 2575 -4885 2615 -4875
rect 2575 -4905 2585 -4885
rect 2605 -4905 2615 -4885
rect 2575 -4915 2615 -4905
rect 2535 -7290 2575 -7280
rect 2535 -7310 2545 -7290
rect 2565 -7310 2575 -7290
rect 2535 -7320 2575 -7310
rect 2600 -7325 2615 -4915
rect 2645 -5785 2685 -5775
rect 2645 -5805 2655 -5785
rect 2675 -5805 2685 -5785
rect 2645 -5815 2685 -5805
rect 2600 -7335 2640 -7325
rect 2600 -7355 2610 -7335
rect 2630 -7355 2640 -7335
rect 2600 -7365 2640 -7355
rect 2670 -7370 2685 -5815
rect 2740 -6525 2780 -6515
rect 2740 -6545 2750 -6525
rect 2770 -6545 2780 -6525
rect 2740 -6555 2780 -6545
rect 2670 -7380 2710 -7370
rect 2670 -7400 2680 -7380
rect 2700 -7400 2710 -7380
rect 2670 -7410 2710 -7400
rect 2740 -7420 2755 -6555
rect 6210 -6675 6225 -665
rect 6825 -1050 6840 -370
rect 30425 -1115 30440 1315
rect 32890 1340 32930 1350
rect 32890 1320 32900 1340
rect 32920 1320 32930 1340
rect 32890 1310 32930 1320
rect 30575 435 30590 740
rect 30550 425 30590 435
rect 30550 405 30560 425
rect 30580 405 30590 425
rect 30550 395 30590 405
rect 32915 -1090 32930 1310
rect 35380 1335 35420 1345
rect 35380 1315 35390 1335
rect 35410 1315 35420 1335
rect 35380 1305 35420 1315
rect 37870 1335 37910 1345
rect 37870 1315 37880 1335
rect 37900 1315 37910 1335
rect 37870 1305 37910 1315
rect 40360 1335 40400 1345
rect 40360 1315 40370 1335
rect 40390 1315 40400 1335
rect 40360 1305 40400 1315
rect 42850 1335 42890 1345
rect 42850 1315 42860 1335
rect 42880 1315 42890 1335
rect 42850 1305 42890 1315
rect 45340 1335 45380 1345
rect 45340 1315 45350 1335
rect 45370 1315 45380 1335
rect 45340 1305 45380 1315
rect 33065 435 33080 735
rect 33040 425 33080 435
rect 33040 405 33050 425
rect 33070 405 33080 425
rect 33040 395 33080 405
rect 35405 -1050 35420 1305
rect 35555 435 35570 735
rect 35530 425 35570 435
rect 35530 405 35540 425
rect 35560 405 35570 425
rect 35530 395 35570 405
rect 37895 -1010 37910 1305
rect 38045 435 38060 735
rect 38020 425 38060 435
rect 38020 405 38030 425
rect 38050 405 38060 425
rect 38020 395 38060 405
rect 40385 -970 40400 1305
rect 40535 435 40550 735
rect 40510 425 40550 435
rect 40510 405 40520 425
rect 40540 405 40550 425
rect 40510 395 40550 405
rect 42875 -930 42890 1305
rect 43025 435 43040 735
rect 43000 425 43040 435
rect 43000 405 43010 425
rect 43030 405 43040 425
rect 43000 395 43040 405
rect 45365 -890 45380 1305
rect 46790 945 46830 955
rect 46790 925 46800 945
rect 46820 925 46830 945
rect 46790 915 46830 925
rect 46790 856 46810 915
rect 46143 835 46810 856
rect 46143 833 46806 835
rect 45515 435 45530 735
rect 45490 425 45530 435
rect 45490 405 45500 425
rect 45520 405 45530 425
rect 45490 395 45530 405
rect 46143 364 46166 833
rect 45535 345 46166 364
rect 45535 -35 45554 345
rect 46143 343 46166 345
rect 7845 -1125 7885 -1115
rect 7845 -1145 7855 -1125
rect 7875 -1140 7885 -1125
rect 28070 -1130 30440 -1115
rect 30560 -1105 32930 -1090
rect 33050 -1065 35420 -1050
rect 35540 -1025 37910 -1010
rect 38030 -985 40400 -970
rect 40520 -945 42890 -930
rect 43010 -905 45380 -890
rect 45500 -54 45554 -35
rect 7875 -1145 8010 -1140
rect 7845 -1155 8010 -1145
rect 6185 -6685 6225 -6675
rect 6185 -6705 6195 -6685
rect 6215 -6705 6225 -6685
rect 6185 -6715 6225 -6705
rect 6250 -1285 6290 -1275
rect 6250 -1305 6260 -1285
rect 6280 -1305 6290 -1285
rect 6250 -1315 6290 -1305
rect 6250 -6740 6265 -1315
rect 6310 -2185 6350 -2175
rect 6310 -2205 6320 -2185
rect 6340 -2205 6350 -2185
rect 6310 -2215 6350 -2205
rect 6225 -6750 6265 -6740
rect 6225 -6770 6235 -6750
rect 6255 -6770 6265 -6750
rect 6225 -6780 6265 -6770
rect 6335 -6800 6350 -2215
rect 6380 -3085 6420 -3075
rect 6380 -3105 6390 -3085
rect 6410 -3105 6420 -3085
rect 6380 -3115 6420 -3105
rect 6335 -6810 6375 -6800
rect 6335 -6830 6345 -6810
rect 6365 -6830 6375 -6810
rect 6335 -6840 6375 -6830
rect 6405 -6845 6420 -3115
rect 6445 -3985 6485 -3975
rect 6445 -4005 6455 -3985
rect 6475 -4005 6485 -3985
rect 6445 -4015 6485 -4005
rect 6405 -6855 6445 -6845
rect 6405 -6875 6415 -6855
rect 6435 -6875 6445 -6855
rect 6405 -6885 6445 -6875
rect 6470 -6890 6485 -4015
rect 6510 -4885 6550 -4875
rect 6510 -4905 6520 -4885
rect 6540 -4905 6550 -4885
rect 6510 -4915 6550 -4905
rect 6470 -6900 6510 -6890
rect 6470 -6920 6480 -6900
rect 6500 -6920 6510 -6900
rect 6470 -6930 6510 -6920
rect 6535 -6935 6550 -4915
rect 7995 -4985 8010 -1155
rect 8040 -1285 8080 -1275
rect 8040 -1305 8050 -1285
rect 8070 -1305 8080 -1285
rect 8040 -1315 8080 -1305
rect 8040 -4760 8055 -1315
rect 28070 -1350 28085 -1130
rect 30560 -1355 30575 -1105
rect 33050 -1360 33065 -1065
rect 35540 -1360 35555 -1025
rect 38030 -1360 38045 -985
rect 40520 -1360 40535 -945
rect 43010 -1360 43025 -905
rect 45500 -1360 45515 -54
rect 8085 -2185 8125 -2175
rect 8085 -2205 8095 -2185
rect 8115 -2205 8125 -2185
rect 8085 -2215 8125 -2205
rect 8085 -4720 8100 -2215
rect 8135 -3085 8175 -3075
rect 8135 -3105 8145 -3085
rect 8165 -3105 8175 -3085
rect 8135 -3115 8175 -3105
rect 28085 -3110 28100 -2755
rect 30575 -3065 30590 -2760
rect 33065 -3065 33080 -2765
rect 35555 -3065 35570 -2765
rect 38045 -3065 38060 -2765
rect 40535 -3065 40550 -2765
rect 43025 -3065 43040 -2765
rect 45515 -3065 45530 -2765
rect 30550 -3075 30590 -3065
rect 30550 -3095 30560 -3075
rect 30580 -3095 30590 -3075
rect 30550 -3105 30590 -3095
rect 33040 -3075 33080 -3065
rect 33040 -3095 33050 -3075
rect 33070 -3095 33080 -3075
rect 33040 -3105 33080 -3095
rect 35530 -3075 35570 -3065
rect 35530 -3095 35540 -3075
rect 35560 -3095 35570 -3075
rect 35530 -3105 35570 -3095
rect 38020 -3075 38060 -3065
rect 38020 -3095 38030 -3075
rect 38050 -3095 38060 -3075
rect 38020 -3105 38060 -3095
rect 40510 -3075 40550 -3065
rect 40510 -3095 40520 -3075
rect 40540 -3095 40550 -3075
rect 40510 -3105 40550 -3095
rect 43000 -3075 43040 -3065
rect 43000 -3095 43010 -3075
rect 43030 -3095 43040 -3075
rect 43000 -3105 43040 -3095
rect 45490 -3075 45530 -3065
rect 45490 -3095 45500 -3075
rect 45520 -3095 45530 -3075
rect 45490 -3105 45530 -3095
rect 8135 -4680 8150 -3115
rect 28060 -3120 28100 -3110
rect 28060 -3140 28070 -3120
rect 28090 -3140 28100 -3120
rect 28060 -3150 28100 -3140
rect 8185 -3985 8225 -3975
rect 8185 -4005 8195 -3985
rect 8215 -4005 8225 -3985
rect 8185 -4015 8225 -4005
rect 8185 -4640 8200 -4015
rect 25915 -4020 25955 -4010
rect 25915 -4040 25925 -4020
rect 25945 -4040 25955 -4020
rect 25915 -4050 25955 -4040
rect 8375 -4505 8415 -4495
rect 8375 -4525 8385 -4505
rect 8405 -4520 8415 -4505
rect 8405 -4525 25440 -4520
rect 8375 -4535 25440 -4525
rect 8310 -4545 8350 -4535
rect 8310 -4565 8320 -4545
rect 8340 -4560 8350 -4545
rect 8340 -4565 22950 -4560
rect 8310 -4575 22950 -4565
rect 8245 -4585 8285 -4575
rect 8245 -4605 8255 -4585
rect 8275 -4600 8285 -4585
rect 8275 -4605 20460 -4600
rect 8245 -4615 20460 -4605
rect 8185 -4655 17970 -4640
rect 8135 -4695 15480 -4680
rect 8085 -4735 12990 -4720
rect 8040 -4775 10500 -4760
rect 10485 -4990 10500 -4775
rect 12975 -4995 12990 -4735
rect 15465 -4995 15480 -4695
rect 17955 -4995 17970 -4655
rect 20445 -4995 20460 -4615
rect 22935 -4995 22950 -4575
rect 25425 -4995 25440 -4535
rect 25915 -4805 25930 -4050
rect 25980 -4070 26020 -4060
rect 25980 -4090 25990 -4070
rect 26010 -4090 26020 -4070
rect 25980 -4100 26020 -4090
rect 25980 -4760 25995 -4100
rect 26050 -4115 26090 -4105
rect 26050 -4135 26060 -4115
rect 26080 -4135 26090 -4115
rect 26050 -4145 26090 -4135
rect 26050 -4720 26065 -4145
rect 26130 -4165 26170 -4155
rect 26130 -4185 26140 -4165
rect 26160 -4185 26170 -4165
rect 26130 -4195 26170 -4185
rect 26130 -4680 26145 -4195
rect 26195 -4215 26235 -4205
rect 26195 -4235 26205 -4215
rect 26225 -4235 26235 -4215
rect 26195 -4245 26235 -4235
rect 26195 -4640 26210 -4245
rect 26265 -4260 26305 -4250
rect 26265 -4280 26275 -4260
rect 26295 -4280 26305 -4260
rect 26265 -4290 26305 -4280
rect 26265 -4600 26280 -4290
rect 26335 -4305 26375 -4295
rect 26335 -4325 26345 -4305
rect 26365 -4325 26375 -4305
rect 26335 -4335 26375 -4325
rect 26335 -4560 26350 -4335
rect 27860 -4505 27900 -4495
rect 27860 -4525 27870 -4505
rect 27890 -4520 27900 -4505
rect 27890 -4525 45515 -4520
rect 27860 -4535 45515 -4525
rect 26335 -4575 43025 -4560
rect 26265 -4615 40535 -4600
rect 26195 -4655 38045 -4640
rect 26130 -4695 35555 -4680
rect 26050 -4735 33065 -4720
rect 25980 -4775 30575 -4760
rect 25915 -4820 28085 -4805
rect 28070 -4980 28085 -4820
rect 30560 -4985 30575 -4775
rect 33050 -4990 33065 -4735
rect 35540 -4990 35555 -4695
rect 38030 -4990 38045 -4655
rect 40520 -4990 40535 -4615
rect 43010 -4990 43025 -4575
rect 45500 -4990 45515 -4535
rect 6580 -5785 6620 -5775
rect 6580 -5805 6590 -5785
rect 6610 -5805 6620 -5785
rect 6580 -5815 6620 -5805
rect 6535 -6945 6575 -6935
rect 6535 -6965 6545 -6945
rect 6565 -6965 6575 -6945
rect 6535 -6975 6575 -6965
rect 6605 -6980 6620 -5815
rect 6675 -6545 6715 -6535
rect 6675 -6565 6685 -6545
rect 6705 -6565 6715 -6545
rect 6675 -6575 6715 -6565
rect 6605 -6990 6645 -6980
rect 6605 -7010 6615 -6990
rect 6635 -7010 6645 -6990
rect 6605 -7020 6645 -7010
rect 6675 -7025 6690 -6575
rect 8010 -6695 8025 -6390
rect 10500 -6695 10515 -6395
rect 12990 -6695 13005 -6400
rect 15480 -6695 15495 -6400
rect 17970 -6695 17985 -6400
rect 20460 -6695 20475 -6400
rect 22950 -6695 22965 -6400
rect 25440 -6695 25455 -6400
rect 7985 -6705 8025 -6695
rect 7985 -6725 7995 -6705
rect 8015 -6725 8025 -6705
rect 7985 -6735 8025 -6725
rect 10475 -6705 10515 -6695
rect 10475 -6725 10485 -6705
rect 10505 -6725 10515 -6705
rect 10475 -6735 10515 -6725
rect 12965 -6705 13005 -6695
rect 12965 -6725 12975 -6705
rect 12995 -6725 13005 -6705
rect 12965 -6735 13005 -6725
rect 15455 -6705 15495 -6695
rect 15455 -6725 15465 -6705
rect 15485 -6725 15495 -6705
rect 15455 -6735 15495 -6725
rect 17945 -6705 17985 -6695
rect 17945 -6725 17955 -6705
rect 17975 -6725 17985 -6705
rect 17945 -6735 17985 -6725
rect 20435 -6705 20475 -6695
rect 20435 -6725 20445 -6705
rect 20465 -6725 20475 -6705
rect 20435 -6735 20475 -6725
rect 22925 -6705 22965 -6695
rect 22925 -6725 22935 -6705
rect 22955 -6725 22965 -6705
rect 22925 -6735 22965 -6725
rect 25415 -6705 25455 -6695
rect 25415 -6725 25425 -6705
rect 25445 -6725 25455 -6705
rect 25415 -6735 25455 -6725
rect 28085 -6740 28100 -6385
rect 30575 -6695 30590 -6390
rect 33065 -6695 33080 -6395
rect 35555 -6695 35570 -6395
rect 38045 -6695 38060 -6395
rect 40535 -6695 40550 -6395
rect 43025 -6695 43040 -6395
rect 45515 -6695 45530 -6395
rect 30550 -6705 30590 -6695
rect 30550 -6725 30560 -6705
rect 30580 -6725 30590 -6705
rect 30550 -6735 30590 -6725
rect 33040 -6705 33080 -6695
rect 33040 -6725 33050 -6705
rect 33070 -6725 33080 -6705
rect 33040 -6735 33080 -6725
rect 35530 -6705 35570 -6695
rect 35530 -6725 35540 -6705
rect 35560 -6725 35570 -6705
rect 35530 -6735 35570 -6725
rect 38020 -6705 38060 -6695
rect 38020 -6725 38030 -6705
rect 38050 -6725 38060 -6705
rect 38020 -6735 38060 -6725
rect 40510 -6705 40550 -6695
rect 40510 -6725 40520 -6705
rect 40540 -6725 40550 -6705
rect 40510 -6735 40550 -6725
rect 43000 -6705 43040 -6695
rect 43000 -6725 43010 -6705
rect 43030 -6725 43040 -6705
rect 43000 -6735 43040 -6725
rect 45490 -6705 45530 -6695
rect 45490 -6725 45500 -6705
rect 45520 -6725 45530 -6705
rect 45490 -6735 45530 -6725
rect 28060 -6750 28100 -6740
rect 28060 -6770 28070 -6750
rect 28090 -6770 28100 -6750
rect 28060 -6780 28100 -6770
rect 6675 -7035 6715 -7025
rect 6675 -7055 6685 -7035
rect 6705 -7055 6715 -7035
rect 6675 -7065 6715 -7055
rect 2740 -7430 2780 -7420
rect 2740 -7450 2750 -7430
rect 2770 -7450 2780 -7430
rect 2740 -7460 2780 -7450
rect 125 -7480 165 -7470
rect 125 -7500 135 -7480
rect 155 -7500 165 -7480
rect 125 -7510 165 -7500
rect 1255 -7480 1295 -7470
rect 1255 -7500 1265 -7480
rect 1285 -7500 1295 -7480
rect 1255 -7510 1295 -7500
rect 2935 -7480 2975 -7470
rect 2935 -7500 2945 -7480
rect 2965 -7500 2975 -7480
rect 2935 -7510 2975 -7500
rect 4065 -7480 4105 -7470
rect 4065 -7500 4075 -7480
rect 4095 -7500 4105 -7480
rect 4065 -7510 4105 -7500
rect 5170 -7480 5210 -7470
rect 5170 -7500 5180 -7480
rect 5200 -7500 5210 -7480
rect 5170 -7510 5210 -7500
rect 125 -8180 140 -7510
rect 1255 -8180 1270 -7510
rect 2250 -7775 2290 -7765
rect 2250 -7795 2260 -7775
rect 2280 -7795 2290 -7775
rect 2250 -7805 2290 -7795
rect 2275 -14205 2290 -7805
rect 2935 -8180 2950 -7510
rect 4065 -8180 4080 -7510
rect 5195 -8180 5210 -7510
rect 6825 -7480 6865 -7470
rect 6825 -7500 6835 -7480
rect 6855 -7500 6865 -7480
rect 6825 -7510 6865 -7500
rect 6185 -7775 6225 -7765
rect 6185 -7795 6195 -7775
rect 6215 -7795 6225 -7775
rect 6185 -7805 6225 -7795
rect 2250 -14215 2290 -14205
rect 2250 -14235 2260 -14215
rect 2280 -14235 2290 -14215
rect 2250 -14245 2290 -14235
rect 2315 -8425 2355 -8415
rect 2315 -8445 2325 -8425
rect 2345 -8445 2355 -8425
rect 2315 -8455 2355 -8445
rect 2315 -14270 2330 -8455
rect 2375 -9325 2415 -9315
rect 2375 -9345 2385 -9325
rect 2405 -9345 2415 -9325
rect 2375 -9355 2415 -9345
rect 2290 -14280 2330 -14270
rect 2290 -14300 2300 -14280
rect 2320 -14300 2330 -14280
rect 2290 -14310 2330 -14300
rect 2400 -14330 2415 -9355
rect 2445 -10225 2485 -10215
rect 2445 -10245 2455 -10225
rect 2475 -10245 2485 -10225
rect 2445 -10255 2485 -10245
rect 2400 -14340 2440 -14330
rect 2400 -14360 2410 -14340
rect 2430 -14360 2440 -14340
rect 2400 -14370 2440 -14360
rect 2470 -14375 2485 -10255
rect 2510 -11125 2550 -11115
rect 2510 -11145 2520 -11125
rect 2540 -11145 2550 -11125
rect 2510 -11155 2550 -11145
rect 2470 -14385 2510 -14375
rect 2470 -14405 2480 -14385
rect 2500 -14405 2510 -14385
rect 2470 -14415 2510 -14405
rect 2535 -14420 2550 -11155
rect 2575 -12025 2615 -12015
rect 2575 -12045 2585 -12025
rect 2605 -12045 2615 -12025
rect 2575 -12055 2615 -12045
rect 2535 -14430 2575 -14420
rect 2535 -14450 2545 -14430
rect 2565 -14450 2575 -14430
rect 2535 -14460 2575 -14450
rect 2600 -14465 2615 -12055
rect 2645 -12925 2685 -12915
rect 2645 -12945 2655 -12925
rect 2675 -12945 2685 -12925
rect 2645 -12955 2685 -12945
rect 2600 -14475 2640 -14465
rect 2600 -14495 2610 -14475
rect 2630 -14495 2640 -14475
rect 2600 -14505 2640 -14495
rect 2670 -14510 2685 -12955
rect 2740 -13665 2780 -13655
rect 2740 -13685 2750 -13665
rect 2770 -13685 2780 -13665
rect 2740 -13695 2780 -13685
rect 2670 -14520 2710 -14510
rect 2670 -14540 2680 -14520
rect 2700 -14540 2710 -14520
rect 2670 -14550 2710 -14540
rect 2740 -14560 2755 -13695
rect 6210 -13815 6225 -7805
rect 6825 -8190 6840 -7510
rect 30345 -8225 30385 -8215
rect 30345 -8245 30355 -8225
rect 30375 -8245 30385 -8225
rect 30345 -8255 30385 -8245
rect 32835 -8225 32875 -8215
rect 32835 -8245 32845 -8225
rect 32865 -8245 32875 -8225
rect 32835 -8255 32875 -8245
rect 35325 -8225 35365 -8215
rect 35325 -8245 35335 -8225
rect 35355 -8245 35365 -8225
rect 35325 -8255 35365 -8245
rect 37815 -8225 37855 -8215
rect 37815 -8245 37825 -8225
rect 37845 -8245 37855 -8225
rect 37815 -8255 37855 -8245
rect 40305 -8225 40345 -8215
rect 40305 -8245 40315 -8225
rect 40335 -8245 40345 -8225
rect 40305 -8255 40345 -8245
rect 42795 -8225 42835 -8215
rect 42795 -8245 42805 -8225
rect 42825 -8245 42835 -8225
rect 42795 -8255 42835 -8245
rect 45285 -8225 45325 -8215
rect 45285 -8245 45295 -8225
rect 45315 -8245 45325 -8225
rect 45285 -8255 45325 -8245
rect 47775 -8225 47815 -8215
rect 47775 -8245 47785 -8225
rect 47805 -8245 47815 -8225
rect 47775 -8255 47815 -8245
rect 7845 -8265 7885 -8255
rect 7845 -8285 7855 -8265
rect 7875 -8280 7885 -8265
rect 7875 -8285 8010 -8280
rect 7845 -8295 8010 -8285
rect 6185 -13825 6225 -13815
rect 6185 -13845 6195 -13825
rect 6215 -13845 6225 -13825
rect 6185 -13855 6225 -13845
rect 6250 -8425 6290 -8415
rect 6250 -8445 6260 -8425
rect 6280 -8445 6290 -8425
rect 6250 -8455 6290 -8445
rect 6250 -13880 6265 -8455
rect 6310 -9325 6350 -9315
rect 6310 -9345 6320 -9325
rect 6340 -9345 6350 -9325
rect 6310 -9355 6350 -9345
rect 6225 -13890 6265 -13880
rect 6225 -13910 6235 -13890
rect 6255 -13910 6265 -13890
rect 6225 -13920 6265 -13910
rect 6335 -13940 6350 -9355
rect 6380 -10225 6420 -10215
rect 6380 -10245 6390 -10225
rect 6410 -10245 6420 -10225
rect 6380 -10255 6420 -10245
rect 6335 -13950 6375 -13940
rect 6335 -13970 6345 -13950
rect 6365 -13970 6375 -13950
rect 6335 -13980 6375 -13970
rect 6405 -13985 6420 -10255
rect 6445 -11125 6485 -11115
rect 6445 -11145 6455 -11125
rect 6475 -11145 6485 -11125
rect 6445 -11155 6485 -11145
rect 6405 -13995 6445 -13985
rect 6405 -14015 6415 -13995
rect 6435 -14015 6445 -13995
rect 6405 -14025 6445 -14015
rect 6470 -14030 6485 -11155
rect 6510 -12025 6550 -12015
rect 6510 -12045 6520 -12025
rect 6540 -12045 6550 -12025
rect 6510 -12055 6550 -12045
rect 6470 -14040 6510 -14030
rect 6470 -14060 6480 -14040
rect 6500 -14060 6510 -14040
rect 6470 -14070 6510 -14060
rect 6535 -14075 6550 -12055
rect 7995 -12125 8010 -8295
rect 8040 -8425 8080 -8415
rect 8040 -8445 8050 -8425
rect 8070 -8445 8080 -8425
rect 8040 -8455 8080 -8445
rect 8040 -11900 8055 -8455
rect 30355 -8650 30370 -8255
rect 32845 -8610 32860 -8255
rect 35335 -8570 35350 -8255
rect 37825 -8530 37840 -8255
rect 40315 -8490 40330 -8255
rect 42805 -8450 42820 -8255
rect 45295 -8410 45310 -8255
rect 47785 -8400 47800 -8255
rect 28070 -8665 30370 -8650
rect 30560 -8625 32860 -8610
rect 33050 -8585 35350 -8570
rect 35540 -8545 37840 -8530
rect 38030 -8505 40330 -8490
rect 40520 -8465 42820 -8450
rect 43010 -8425 45310 -8410
rect 45500 -8415 47800 -8400
rect 28070 -8870 28085 -8665
rect 30560 -8875 30575 -8625
rect 33050 -8880 33065 -8585
rect 35540 -8880 35555 -8545
rect 38030 -8880 38045 -8505
rect 40520 -8880 40535 -8465
rect 43010 -8880 43025 -8425
rect 45500 -8880 45515 -8415
rect 8085 -9325 8125 -9315
rect 8085 -9345 8095 -9325
rect 8115 -9345 8125 -9325
rect 8085 -9355 8125 -9345
rect 8085 -11860 8100 -9355
rect 8135 -10225 8175 -10215
rect 8135 -10245 8145 -10225
rect 8165 -10245 8175 -10225
rect 8135 -10255 8175 -10245
rect 8135 -11820 8150 -10255
rect 28085 -10630 28100 -10275
rect 30575 -10585 30590 -10280
rect 33065 -10585 33080 -10285
rect 35555 -10585 35570 -10285
rect 38045 -10585 38060 -10285
rect 40535 -10585 40550 -10285
rect 43025 -10585 43040 -10285
rect 45515 -10585 45530 -10285
rect 30550 -10595 30590 -10585
rect 30550 -10615 30560 -10595
rect 30580 -10615 30590 -10595
rect 30550 -10625 30590 -10615
rect 33040 -10595 33080 -10585
rect 33040 -10615 33050 -10595
rect 33070 -10615 33080 -10595
rect 33040 -10625 33080 -10615
rect 35530 -10595 35570 -10585
rect 35530 -10615 35540 -10595
rect 35560 -10615 35570 -10595
rect 35530 -10625 35570 -10615
rect 38020 -10595 38060 -10585
rect 38020 -10615 38030 -10595
rect 38050 -10615 38060 -10595
rect 38020 -10625 38060 -10615
rect 40510 -10595 40550 -10585
rect 40510 -10615 40520 -10595
rect 40540 -10615 40550 -10595
rect 40510 -10625 40550 -10615
rect 43000 -10595 43040 -10585
rect 43000 -10615 43010 -10595
rect 43030 -10615 43040 -10595
rect 43000 -10625 43040 -10615
rect 45490 -10595 45530 -10585
rect 45490 -10615 45500 -10595
rect 45520 -10615 45530 -10595
rect 45490 -10625 45530 -10615
rect 28060 -10640 28100 -10630
rect 28060 -10660 28070 -10640
rect 28090 -10660 28100 -10640
rect 28060 -10670 28100 -10660
rect 8185 -11125 8225 -11115
rect 8185 -11145 8195 -11125
rect 8215 -11145 8225 -11125
rect 8185 -11155 8225 -11145
rect 8185 -11780 8200 -11155
rect 25915 -11160 25955 -11150
rect 25915 -11180 25925 -11160
rect 25945 -11180 25955 -11160
rect 25915 -11190 25955 -11180
rect 8375 -11645 8415 -11635
rect 8375 -11665 8385 -11645
rect 8405 -11660 8415 -11645
rect 8405 -11665 25440 -11660
rect 8375 -11675 25440 -11665
rect 8310 -11685 8350 -11675
rect 8310 -11705 8320 -11685
rect 8340 -11700 8350 -11685
rect 8340 -11705 22950 -11700
rect 8310 -11715 22950 -11705
rect 8245 -11725 8285 -11715
rect 8245 -11745 8255 -11725
rect 8275 -11740 8285 -11725
rect 8275 -11745 20460 -11740
rect 8245 -11755 20460 -11745
rect 8185 -11795 17970 -11780
rect 8135 -11835 15480 -11820
rect 8085 -11875 12990 -11860
rect 8040 -11915 10500 -11900
rect 10485 -12130 10500 -11915
rect 12975 -12135 12990 -11875
rect 15465 -12135 15480 -11835
rect 17955 -12135 17970 -11795
rect 20445 -12135 20460 -11755
rect 22935 -12135 22950 -11715
rect 25425 -12135 25440 -11675
rect 25915 -11945 25930 -11190
rect 25980 -11210 26020 -11200
rect 25980 -11230 25990 -11210
rect 26010 -11230 26020 -11210
rect 25980 -11240 26020 -11230
rect 25980 -11900 25995 -11240
rect 26050 -11255 26090 -11245
rect 26050 -11275 26060 -11255
rect 26080 -11275 26090 -11255
rect 26050 -11285 26090 -11275
rect 26050 -11860 26065 -11285
rect 26130 -11305 26170 -11295
rect 26130 -11325 26140 -11305
rect 26160 -11325 26170 -11305
rect 26130 -11335 26170 -11325
rect 26130 -11820 26145 -11335
rect 26195 -11355 26235 -11345
rect 26195 -11375 26205 -11355
rect 26225 -11375 26235 -11355
rect 26195 -11385 26235 -11375
rect 26195 -11780 26210 -11385
rect 26265 -11400 26305 -11390
rect 26265 -11420 26275 -11400
rect 26295 -11420 26305 -11400
rect 26265 -11430 26305 -11420
rect 26265 -11740 26280 -11430
rect 26335 -11445 26375 -11435
rect 26335 -11465 26345 -11445
rect 26365 -11465 26375 -11445
rect 26335 -11475 26375 -11465
rect 26335 -11700 26350 -11475
rect 27860 -11645 27900 -11635
rect 27860 -11665 27870 -11645
rect 27890 -11660 27900 -11645
rect 27890 -11665 45515 -11660
rect 27860 -11675 45515 -11665
rect 26335 -11715 43025 -11700
rect 26265 -11755 40535 -11740
rect 26195 -11795 38045 -11780
rect 26130 -11835 35555 -11820
rect 26050 -11875 33065 -11860
rect 25980 -11915 30575 -11900
rect 25915 -11960 28085 -11945
rect 28070 -12120 28085 -11960
rect 30560 -12125 30575 -11915
rect 33050 -12130 33065 -11875
rect 35540 -12130 35555 -11835
rect 38030 -12130 38045 -11795
rect 40520 -12130 40535 -11755
rect 43010 -12130 43025 -11715
rect 45500 -12130 45515 -11675
rect 6580 -12925 6620 -12915
rect 6580 -12945 6590 -12925
rect 6610 -12945 6620 -12925
rect 6580 -12955 6620 -12945
rect 6535 -14085 6575 -14075
rect 6535 -14105 6545 -14085
rect 6565 -14105 6575 -14085
rect 6535 -14115 6575 -14105
rect 6605 -14120 6620 -12955
rect 6675 -13685 6715 -13675
rect 6675 -13705 6685 -13685
rect 6705 -13705 6715 -13685
rect 6675 -13715 6715 -13705
rect 6605 -14130 6645 -14120
rect 6605 -14150 6615 -14130
rect 6635 -14150 6645 -14130
rect 6605 -14160 6645 -14150
rect 6675 -14165 6690 -13715
rect 8010 -13835 8025 -13530
rect 10500 -13835 10515 -13535
rect 12990 -13835 13005 -13540
rect 15480 -13835 15495 -13540
rect 17970 -13835 17985 -13540
rect 20460 -13835 20475 -13540
rect 22950 -13835 22965 -13540
rect 25440 -13835 25455 -13540
rect 7985 -13845 8025 -13835
rect 7985 -13865 7995 -13845
rect 8015 -13865 8025 -13845
rect 7985 -13875 8025 -13865
rect 10475 -13845 10515 -13835
rect 10475 -13865 10485 -13845
rect 10505 -13865 10515 -13845
rect 10475 -13875 10515 -13865
rect 12965 -13845 13005 -13835
rect 12965 -13865 12975 -13845
rect 12995 -13865 13005 -13845
rect 12965 -13875 13005 -13865
rect 15455 -13845 15495 -13835
rect 15455 -13865 15465 -13845
rect 15485 -13865 15495 -13845
rect 15455 -13875 15495 -13865
rect 17945 -13845 17985 -13835
rect 17945 -13865 17955 -13845
rect 17975 -13865 17985 -13845
rect 17945 -13875 17985 -13865
rect 20435 -13845 20475 -13835
rect 20435 -13865 20445 -13845
rect 20465 -13865 20475 -13845
rect 20435 -13875 20475 -13865
rect 22925 -13845 22965 -13835
rect 22925 -13865 22935 -13845
rect 22955 -13865 22965 -13845
rect 22925 -13875 22965 -13865
rect 25415 -13845 25455 -13835
rect 25415 -13865 25425 -13845
rect 25445 -13865 25455 -13845
rect 25415 -13875 25455 -13865
rect 28085 -13880 28100 -13525
rect 30575 -13835 30590 -13530
rect 33065 -13835 33080 -13535
rect 35555 -13835 35570 -13535
rect 38045 -13835 38060 -13535
rect 40535 -13835 40550 -13535
rect 43025 -13835 43040 -13535
rect 45515 -13835 45530 -13535
rect 30550 -13845 30590 -13835
rect 30550 -13865 30560 -13845
rect 30580 -13865 30590 -13845
rect 30550 -13875 30590 -13865
rect 33040 -13845 33080 -13835
rect 33040 -13865 33050 -13845
rect 33070 -13865 33080 -13845
rect 33040 -13875 33080 -13865
rect 35530 -13845 35570 -13835
rect 35530 -13865 35540 -13845
rect 35560 -13865 35570 -13845
rect 35530 -13875 35570 -13865
rect 38020 -13845 38060 -13835
rect 38020 -13865 38030 -13845
rect 38050 -13865 38060 -13845
rect 38020 -13875 38060 -13865
rect 40510 -13845 40550 -13835
rect 40510 -13865 40520 -13845
rect 40540 -13865 40550 -13845
rect 40510 -13875 40550 -13865
rect 43000 -13845 43040 -13835
rect 43000 -13865 43010 -13845
rect 43030 -13865 43040 -13845
rect 43000 -13875 43040 -13865
rect 45490 -13845 45530 -13835
rect 45490 -13865 45500 -13845
rect 45520 -13865 45530 -13845
rect 45490 -13875 45530 -13865
rect 28060 -13890 28100 -13880
rect 28060 -13910 28070 -13890
rect 28090 -13910 28100 -13890
rect 28060 -13920 28100 -13910
rect 6675 -14175 6715 -14165
rect 6675 -14195 6685 -14175
rect 6705 -14195 6715 -14175
rect 6675 -14205 6715 -14195
rect 2740 -14570 2780 -14560
rect 2740 -14590 2750 -14570
rect 2770 -14590 2780 -14570
rect 2740 -14600 2780 -14590
<< polycont >>
rect 135 6770 155 6790
rect 1815 6770 1835 6790
rect 2945 6770 2965 6790
rect 4075 6770 4095 6790
rect 5705 6770 5725 6790
rect 6835 6770 6855 6790
rect 1135 6475 1155 6495
rect 5070 6475 5090 6495
rect 1135 35 1155 55
rect 1200 5825 1220 5845
rect 1260 4925 1280 4945
rect 1175 -30 1195 -10
rect 1330 4025 1350 4045
rect 1285 -90 1305 -70
rect 1395 3125 1415 3145
rect 1355 -135 1375 -115
rect 1460 2225 1480 2245
rect 1420 -180 1440 -160
rect 1530 1325 1550 1345
rect 1485 -225 1505 -205
rect 1625 585 1645 605
rect 1555 -270 1575 -250
rect 7855 5985 7875 6005
rect 5070 425 5090 445
rect 5135 5825 5155 5845
rect 5195 4925 5215 4945
rect 5110 360 5130 380
rect 5265 4025 5285 4045
rect 5220 300 5240 320
rect 5330 3125 5350 3145
rect 5290 255 5310 275
rect 5395 2225 5415 2245
rect 5355 210 5375 230
rect 8050 5825 8070 5845
rect 8095 4925 8115 4945
rect 8145 4025 8165 4045
rect 8195 3125 8215 3145
rect 25925 3090 25945 3110
rect 8385 2605 8405 2625
rect 8320 2565 8340 2585
rect 8255 2525 8275 2545
rect 25990 3040 26010 3060
rect 26060 2995 26080 3015
rect 26140 2945 26160 2965
rect 26205 2895 26225 2915
rect 26275 2850 26295 2870
rect 26345 2805 26365 2825
rect 27870 2605 27890 2625
rect 5465 1325 5485 1345
rect 30410 1325 30430 1345
rect 5420 165 5440 185
rect 5560 565 5580 585
rect 5490 120 5510 140
rect 7995 405 8015 425
rect 10485 405 10505 425
rect 12975 405 12995 425
rect 15465 405 15485 425
rect 17955 405 17975 425
rect 20445 405 20465 425
rect 22935 405 22955 425
rect 25425 405 25445 425
rect 28070 360 28090 380
rect 5560 75 5580 95
rect 1625 -320 1645 -300
rect 135 -360 155 -340
rect 1265 -360 1285 -340
rect 2945 -360 2965 -340
rect 4075 -360 4095 -340
rect 5180 -360 5200 -340
rect 2260 -655 2280 -635
rect 6835 -360 6855 -340
rect 6195 -655 6215 -635
rect 2260 -7095 2280 -7075
rect 2325 -1305 2345 -1285
rect 2385 -2205 2405 -2185
rect 2300 -7160 2320 -7140
rect 2455 -3105 2475 -3085
rect 2410 -7220 2430 -7200
rect 2520 -4005 2540 -3985
rect 2480 -7265 2500 -7245
rect 2585 -4905 2605 -4885
rect 2545 -7310 2565 -7290
rect 2655 -5805 2675 -5785
rect 2610 -7355 2630 -7335
rect 2750 -6545 2770 -6525
rect 2680 -7400 2700 -7380
rect 32900 1320 32920 1340
rect 30560 405 30580 425
rect 35390 1315 35410 1335
rect 37880 1315 37900 1335
rect 40370 1315 40390 1335
rect 42860 1315 42880 1335
rect 45350 1315 45370 1335
rect 33050 405 33070 425
rect 35540 405 35560 425
rect 38030 405 38050 425
rect 40520 405 40540 425
rect 43010 405 43030 425
rect 46800 925 46820 945
rect 45500 405 45520 425
rect 7855 -1145 7875 -1125
rect 6195 -6705 6215 -6685
rect 6260 -1305 6280 -1285
rect 6320 -2205 6340 -2185
rect 6235 -6770 6255 -6750
rect 6390 -3105 6410 -3085
rect 6345 -6830 6365 -6810
rect 6455 -4005 6475 -3985
rect 6415 -6875 6435 -6855
rect 6520 -4905 6540 -4885
rect 6480 -6920 6500 -6900
rect 8050 -1305 8070 -1285
rect 8095 -2205 8115 -2185
rect 8145 -3105 8165 -3085
rect 30560 -3095 30580 -3075
rect 33050 -3095 33070 -3075
rect 35540 -3095 35560 -3075
rect 38030 -3095 38050 -3075
rect 40520 -3095 40540 -3075
rect 43010 -3095 43030 -3075
rect 45500 -3095 45520 -3075
rect 28070 -3140 28090 -3120
rect 8195 -4005 8215 -3985
rect 25925 -4040 25945 -4020
rect 8385 -4525 8405 -4505
rect 8320 -4565 8340 -4545
rect 8255 -4605 8275 -4585
rect 25990 -4090 26010 -4070
rect 26060 -4135 26080 -4115
rect 26140 -4185 26160 -4165
rect 26205 -4235 26225 -4215
rect 26275 -4280 26295 -4260
rect 26345 -4325 26365 -4305
rect 27870 -4525 27890 -4505
rect 6590 -5805 6610 -5785
rect 6545 -6965 6565 -6945
rect 6685 -6565 6705 -6545
rect 6615 -7010 6635 -6990
rect 7995 -6725 8015 -6705
rect 10485 -6725 10505 -6705
rect 12975 -6725 12995 -6705
rect 15465 -6725 15485 -6705
rect 17955 -6725 17975 -6705
rect 20445 -6725 20465 -6705
rect 22935 -6725 22955 -6705
rect 25425 -6725 25445 -6705
rect 30560 -6725 30580 -6705
rect 33050 -6725 33070 -6705
rect 35540 -6725 35560 -6705
rect 38030 -6725 38050 -6705
rect 40520 -6725 40540 -6705
rect 43010 -6725 43030 -6705
rect 45500 -6725 45520 -6705
rect 28070 -6770 28090 -6750
rect 6685 -7055 6705 -7035
rect 2750 -7450 2770 -7430
rect 135 -7500 155 -7480
rect 1265 -7500 1285 -7480
rect 2945 -7500 2965 -7480
rect 4075 -7500 4095 -7480
rect 5180 -7500 5200 -7480
rect 2260 -7795 2280 -7775
rect 6835 -7500 6855 -7480
rect 6195 -7795 6215 -7775
rect 2260 -14235 2280 -14215
rect 2325 -8445 2345 -8425
rect 2385 -9345 2405 -9325
rect 2300 -14300 2320 -14280
rect 2455 -10245 2475 -10225
rect 2410 -14360 2430 -14340
rect 2520 -11145 2540 -11125
rect 2480 -14405 2500 -14385
rect 2585 -12045 2605 -12025
rect 2545 -14450 2565 -14430
rect 2655 -12945 2675 -12925
rect 2610 -14495 2630 -14475
rect 2750 -13685 2770 -13665
rect 2680 -14540 2700 -14520
rect 30355 -8245 30375 -8225
rect 32845 -8245 32865 -8225
rect 35335 -8245 35355 -8225
rect 37825 -8245 37845 -8225
rect 40315 -8245 40335 -8225
rect 42805 -8245 42825 -8225
rect 45295 -8245 45315 -8225
rect 47785 -8245 47805 -8225
rect 7855 -8285 7875 -8265
rect 6195 -13845 6215 -13825
rect 6260 -8445 6280 -8425
rect 6320 -9345 6340 -9325
rect 6235 -13910 6255 -13890
rect 6390 -10245 6410 -10225
rect 6345 -13970 6365 -13950
rect 6455 -11145 6475 -11125
rect 6415 -14015 6435 -13995
rect 6520 -12045 6540 -12025
rect 6480 -14060 6500 -14040
rect 8050 -8445 8070 -8425
rect 8095 -9345 8115 -9325
rect 8145 -10245 8165 -10225
rect 30560 -10615 30580 -10595
rect 33050 -10615 33070 -10595
rect 35540 -10615 35560 -10595
rect 38030 -10615 38050 -10595
rect 40520 -10615 40540 -10595
rect 43010 -10615 43030 -10595
rect 45500 -10615 45520 -10595
rect 28070 -10660 28090 -10640
rect 8195 -11145 8215 -11125
rect 25925 -11180 25945 -11160
rect 8385 -11665 8405 -11645
rect 8320 -11705 8340 -11685
rect 8255 -11745 8275 -11725
rect 25990 -11230 26010 -11210
rect 26060 -11275 26080 -11255
rect 26140 -11325 26160 -11305
rect 26205 -11375 26225 -11355
rect 26275 -11420 26295 -11400
rect 26345 -11465 26365 -11445
rect 27870 -11665 27890 -11645
rect 6590 -12945 6610 -12925
rect 6545 -14105 6565 -14085
rect 6685 -13705 6705 -13685
rect 6615 -14150 6635 -14130
rect 7995 -13865 8015 -13845
rect 10485 -13865 10505 -13845
rect 12975 -13865 12995 -13845
rect 15465 -13865 15485 -13845
rect 17955 -13865 17975 -13845
rect 20445 -13865 20465 -13845
rect 22935 -13865 22955 -13845
rect 25425 -13865 25445 -13845
rect 30560 -13865 30580 -13845
rect 33050 -13865 33070 -13845
rect 35540 -13865 35560 -13845
rect 38030 -13865 38050 -13845
rect 40520 -13865 40540 -13845
rect 43010 -13865 43030 -13845
rect 45500 -13865 45520 -13845
rect 28070 -13910 28090 -13890
rect 6685 -14195 6705 -14175
rect 2750 -14590 2770 -14570
<< locali >>
rect 125 6790 165 6800
rect 125 6770 135 6790
rect 155 6780 165 6790
rect 1805 6790 1845 6800
rect 1805 6780 1815 6790
rect 155 6770 1815 6780
rect 1835 6780 1845 6790
rect 2935 6790 2975 6800
rect 2935 6780 2945 6790
rect 1835 6770 2945 6780
rect 2965 6780 2975 6790
rect 4065 6790 4105 6800
rect 4065 6780 4075 6790
rect 2965 6770 4075 6780
rect 4095 6780 4105 6790
rect 5695 6790 5735 6800
rect 5695 6780 5705 6790
rect 4095 6770 5705 6780
rect 5725 6780 5735 6790
rect 6825 6790 6865 6800
rect 6825 6780 6835 6790
rect 5725 6770 6835 6780
rect 6855 6770 6865 6790
rect 125 6760 6865 6770
rect 55 6720 6775 6740
rect 55 6575 75 6720
rect 1735 6580 1755 6720
rect 2865 6580 2885 6720
rect 3995 6580 4015 6720
rect 5620 6580 5640 6720
rect 6755 6580 6775 6720
rect 3975 6560 3985 6580
rect 1125 6495 1900 6505
rect 1125 6475 1135 6495
rect 1155 6485 1900 6495
rect 2805 6485 3060 6505
rect 3935 6485 4145 6505
rect 5060 6495 5800 6505
rect 1155 6475 1165 6485
rect 1125 6465 1165 6475
rect 1125 5975 1145 6465
rect 2805 5980 2825 6485
rect 3935 5995 3955 6485
rect 5060 6475 5070 6495
rect 5090 6485 5800 6495
rect 6695 6485 6915 6505
rect 5090 6475 5100 6485
rect 5060 6465 5100 6475
rect 5065 6000 5085 6465
rect 3930 5980 3955 5995
rect 5060 5975 5085 6000
rect 6695 5975 6715 6485
rect 7845 6005 7885 6015
rect 7845 5985 7855 6005
rect 7875 5985 7885 6005
rect 7845 5975 7885 5985
rect 1190 5845 1230 5855
rect 1190 5835 1200 5845
rect 1135 5825 1200 5835
rect 1220 5835 1230 5845
rect 5125 5845 5165 5855
rect 5125 5835 5135 5845
rect 1220 5825 1825 5835
rect 1135 5815 1825 5825
rect 2815 5815 2970 5835
rect 3950 5815 4100 5835
rect 5085 5825 5135 5835
rect 5155 5835 5165 5845
rect 8040 5845 8080 5855
rect 8040 5835 8050 5845
rect 5155 5825 5730 5835
rect 5085 5815 5730 5825
rect 6710 5815 6855 5835
rect 7845 5825 8050 5835
rect 8070 5825 8080 5845
rect 7845 5815 8080 5825
rect 1250 4945 1290 4955
rect 1250 4935 1260 4945
rect 1140 4925 1260 4935
rect 1280 4935 1290 4945
rect 5185 4945 5225 4955
rect 5185 4935 5195 4945
rect 1280 4925 1830 4935
rect 1140 4915 1830 4925
rect 2820 4915 2975 4935
rect 3955 4915 4105 4935
rect 5085 4925 5195 4935
rect 5215 4935 5225 4945
rect 8085 4945 8125 4955
rect 8085 4935 8095 4945
rect 5215 4925 5730 4935
rect 5085 4915 5730 4925
rect 6710 4915 6855 4935
rect 7845 4925 8095 4935
rect 8115 4925 8125 4945
rect 7845 4915 8125 4925
rect 1320 4045 1360 4055
rect 1320 4035 1330 4045
rect 1140 4025 1330 4035
rect 1350 4035 1360 4045
rect 5255 4045 5295 4055
rect 5255 4035 5265 4045
rect 1350 4025 1830 4035
rect 1140 4015 1830 4025
rect 2815 4015 2970 4035
rect 3950 4015 4100 4035
rect 5085 4025 5265 4035
rect 5285 4035 5295 4045
rect 8135 4045 8175 4055
rect 8135 4035 8145 4045
rect 5285 4025 5730 4035
rect 5085 4015 5730 4025
rect 6715 4015 6860 4035
rect 7845 4025 8145 4035
rect 8165 4025 8175 4045
rect 7845 4015 8175 4025
rect 1385 3145 1425 3155
rect 1385 3135 1395 3145
rect 1140 3125 1395 3135
rect 1415 3135 1425 3145
rect 5320 3145 5360 3155
rect 5320 3135 5330 3145
rect 1415 3125 1830 3135
rect 1140 3115 1830 3125
rect 2820 3115 2975 3135
rect 3950 3115 4100 3135
rect 5085 3125 5330 3135
rect 5350 3135 5360 3145
rect 8185 3145 8225 3155
rect 8185 3135 8195 3145
rect 5350 3125 5730 3135
rect 5085 3115 5730 3125
rect 6710 3115 6855 3135
rect 7845 3125 8195 3135
rect 8215 3125 8225 3145
rect 7845 3115 8225 3125
rect 25915 3110 25955 3120
rect 25915 3105 25925 3110
rect 25445 3090 25925 3105
rect 25945 3090 25955 3110
rect 25445 3080 25955 3090
rect 25445 2695 25470 3080
rect 25980 3060 26020 3070
rect 25980 3055 25990 3060
rect 10365 2670 25470 2695
rect 25495 3040 25990 3055
rect 26010 3040 26020 3060
rect 25495 3030 26020 3040
rect 8375 2625 8415 2635
rect 8375 2605 8385 2625
rect 8405 2605 8415 2625
rect 8375 2595 8415 2605
rect 8310 2585 8350 2595
rect 8310 2565 8320 2585
rect 8340 2565 8350 2585
rect 8310 2555 8350 2565
rect 8245 2545 8285 2555
rect 8245 2535 8255 2545
rect 7845 2525 8255 2535
rect 8275 2525 8285 2545
rect 7845 2515 8285 2525
rect 1450 2245 1490 2255
rect 1450 2235 1460 2245
rect 1130 2225 1460 2235
rect 1480 2235 1490 2245
rect 5385 2245 5425 2255
rect 5385 2235 5395 2245
rect 1480 2225 1835 2235
rect 1130 2215 1835 2225
rect 2820 2215 2975 2235
rect 3940 2215 4090 2235
rect 5085 2225 5395 2235
rect 5415 2235 5425 2245
rect 5415 2225 5730 2235
rect 5085 2215 5730 2225
rect 6705 2215 6850 2235
rect 7845 2215 7865 2515
rect 8310 2490 8330 2555
rect 7890 2470 8330 2490
rect 1520 1345 1560 1355
rect 1520 1335 1530 1345
rect 1135 1325 1530 1335
rect 1550 1335 1560 1345
rect 5455 1345 5495 1355
rect 5455 1335 5465 1345
rect 1550 1325 1830 1335
rect 1135 1315 1830 1325
rect 2810 1315 2965 1335
rect 3950 1315 4100 1335
rect 5085 1325 5465 1335
rect 5485 1335 5495 1345
rect 7890 1335 7910 2470
rect 8375 2445 8395 2595
rect 5485 1325 5730 1335
rect 5085 1315 5730 1325
rect 6710 1315 6855 1335
rect 7835 1315 7910 1335
rect 7935 2425 8395 2445
rect 7935 1025 7955 2425
rect 9245 2105 9250 2110
rect 10365 2105 10385 2670
rect 25495 2645 25520 3030
rect 26050 3015 26090 3025
rect 26050 3010 26060 3015
rect 12855 2620 25520 2645
rect 25540 2995 26060 3010
rect 26080 2995 26090 3015
rect 25540 2985 26090 2995
rect 12855 2105 12875 2620
rect 25540 2595 25565 2985
rect 26130 2965 26170 2975
rect 26130 2960 26140 2965
rect 15345 2570 25565 2595
rect 25585 2945 26140 2960
rect 26160 2945 26170 2965
rect 25585 2935 26170 2945
rect 15345 2105 15365 2570
rect 25585 2545 25610 2935
rect 26195 2915 26235 2925
rect 26195 2910 26205 2915
rect 17835 2520 25610 2545
rect 25630 2895 26205 2910
rect 26225 2895 26235 2915
rect 25630 2885 26235 2895
rect 17835 2105 17855 2520
rect 25630 2490 25655 2885
rect 26265 2870 26305 2880
rect 26265 2865 26275 2870
rect 20325 2465 25655 2490
rect 25680 2850 26275 2865
rect 26295 2850 26305 2870
rect 25680 2840 26305 2850
rect 25680 2820 25710 2840
rect 26335 2825 26375 2835
rect 26335 2820 26345 2825
rect 20325 2105 20345 2465
rect 25680 2440 25705 2820
rect 22815 2415 25705 2440
rect 25730 2805 26345 2820
rect 26365 2805 26375 2825
rect 25730 2795 26375 2805
rect 22815 2105 22835 2415
rect 25730 2390 25755 2795
rect 25305 2365 25755 2390
rect 27860 2625 27900 2635
rect 27860 2605 27870 2625
rect 27890 2605 27900 2625
rect 27860 2595 27900 2605
rect 25305 2105 25325 2365
rect 9310 2085 9330 2105
rect 10365 2085 10450 2105
rect 12855 2085 12940 2105
rect 15345 2085 15430 2105
rect 17835 2085 17920 2105
rect 20325 2085 20410 2105
rect 22815 2085 22900 2105
rect 25305 2085 25390 2105
rect 9305 2080 9330 2085
rect 9305 2075 9325 2080
rect 9300 1910 9305 1915
rect 9295 1890 9305 1910
rect 10430 1645 10450 2085
rect 12920 1640 12940 2085
rect 15410 1635 15430 2085
rect 17900 1635 17920 2085
rect 20390 1635 20410 2085
rect 22880 1635 22900 2085
rect 25370 1635 25390 2085
rect 27860 1635 27885 2595
rect 29375 2090 29405 2115
rect 30500 1650 30540 1670
rect 30520 1355 30540 1650
rect 30400 1345 30540 1355
rect 33010 1350 33030 1665
rect 35480 1640 35520 1660
rect 37970 1640 38010 1660
rect 40460 1640 40500 1660
rect 42950 1640 42990 1660
rect 45445 1640 45480 1660
rect 30400 1325 30410 1345
rect 30430 1335 30540 1345
rect 32890 1340 33030 1350
rect 35500 1345 35520 1640
rect 37990 1345 38010 1640
rect 40480 1345 40500 1640
rect 42970 1345 42990 1640
rect 45460 1345 45480 1640
rect 47935 1345 47955 1660
rect 30430 1325 30440 1335
rect 30400 1315 30440 1325
rect 32890 1320 32900 1340
rect 32920 1330 33030 1340
rect 35380 1335 35520 1345
rect 32920 1320 32930 1330
rect 32890 1310 32930 1320
rect 35380 1315 35390 1335
rect 35410 1325 35520 1335
rect 37870 1335 38010 1345
rect 35410 1315 35420 1325
rect 35380 1305 35420 1315
rect 37870 1315 37880 1335
rect 37900 1325 38010 1335
rect 40360 1335 40500 1345
rect 37900 1315 37910 1325
rect 37870 1305 37910 1315
rect 40360 1315 40370 1335
rect 40390 1325 40500 1335
rect 42850 1335 42990 1345
rect 40390 1315 40400 1325
rect 40360 1305 40400 1315
rect 42850 1315 42860 1335
rect 42880 1325 42990 1335
rect 45340 1335 45480 1345
rect 42880 1315 42890 1325
rect 42850 1305 42890 1315
rect 45340 1315 45350 1335
rect 45370 1325 45480 1335
rect 46800 1325 47955 1345
rect 45370 1315 45380 1325
rect 45340 1305 45380 1315
rect 1145 1005 1655 1025
rect 1635 615 1655 1005
rect 1615 605 1655 615
rect 1615 585 1625 605
rect 1645 595 1655 605
rect 2800 595 2825 1020
rect 3930 1005 3955 1020
rect 3935 595 3955 1005
rect 5065 595 5085 1015
rect 6695 595 6715 1010
rect 7835 1005 7955 1025
rect 46800 955 46820 1325
rect 46790 945 46830 955
rect 46790 925 46800 945
rect 46820 925 46830 945
rect 46790 915 46830 925
rect 1645 585 1890 595
rect 1615 575 1890 585
rect 2800 575 3020 595
rect 3935 575 4165 595
rect 5065 585 5780 595
rect 5065 575 5560 585
rect 5550 565 5560 575
rect 5580 575 5780 585
rect 6695 575 6920 595
rect 5580 565 5590 575
rect 5550 555 5590 565
rect 5060 445 5100 455
rect 5060 425 5070 445
rect 5090 435 5100 445
rect 5090 425 8025 435
rect 5060 415 7995 425
rect 7985 405 7995 415
rect 8015 415 8025 425
rect 10475 425 10515 435
rect 8015 405 8030 415
rect 7985 395 8030 405
rect 10475 405 10485 425
rect 10505 405 10515 425
rect 10475 395 10515 405
rect 12965 425 13005 435
rect 12965 405 12975 425
rect 12995 405 13005 425
rect 12965 395 13005 405
rect 15455 425 15495 435
rect 15455 405 15465 425
rect 15485 405 15495 425
rect 15455 395 15495 405
rect 17945 425 17985 435
rect 17945 405 17955 425
rect 17975 405 17985 425
rect 17945 395 17985 405
rect 20435 425 20475 435
rect 20435 405 20445 425
rect 20465 405 20475 425
rect 20435 395 20475 405
rect 22925 425 22965 435
rect 22925 405 22935 425
rect 22955 405 22965 425
rect 22925 395 22965 405
rect 25415 425 25455 435
rect 25415 405 25425 425
rect 25445 405 25455 425
rect 25415 395 25455 405
rect 30550 425 30590 435
rect 30550 405 30560 425
rect 30580 415 30590 425
rect 33040 425 33080 435
rect 30580 405 30595 415
rect 30550 395 30595 405
rect 33040 405 33050 425
rect 33070 420 33080 425
rect 35530 425 35570 435
rect 33070 405 33090 420
rect 33040 395 33090 405
rect 35530 405 35540 425
rect 35560 415 35570 425
rect 38020 425 38060 435
rect 35560 405 35575 415
rect 35530 395 35575 405
rect 38020 405 38030 425
rect 38050 415 38060 425
rect 40510 425 40550 435
rect 38050 405 38065 415
rect 38020 395 38065 405
rect 40510 405 40520 425
rect 40540 415 40550 425
rect 43000 425 43040 435
rect 40540 405 40555 415
rect 40510 395 40555 405
rect 43000 405 43010 425
rect 43030 420 43040 425
rect 45490 425 45530 435
rect 43030 405 43045 420
rect 43000 395 43045 405
rect 45490 405 45500 425
rect 45520 415 45530 425
rect 45520 405 45535 415
rect 45490 395 45535 405
rect 5100 380 5140 390
rect 5100 360 5110 380
rect 5130 370 5140 380
rect 10475 370 10495 395
rect 5130 360 10495 370
rect 5100 350 10495 360
rect 12965 330 12990 395
rect 5210 320 12990 330
rect 5210 300 5220 320
rect 5240 310 12990 320
rect 5240 300 5250 310
rect 5210 290 5250 300
rect 15455 285 15475 395
rect 5280 275 15475 285
rect 5280 255 5290 275
rect 5310 265 15475 275
rect 5310 255 5320 265
rect 5280 245 5320 255
rect 17945 240 17965 395
rect 5345 230 17965 240
rect 5345 210 5355 230
rect 5375 220 17965 230
rect 5375 210 5385 220
rect 5345 200 5385 210
rect 20435 195 20455 395
rect 5410 185 20455 195
rect 5410 165 5420 185
rect 5440 175 20455 185
rect 5440 165 5450 175
rect 5410 155 5450 165
rect 22925 150 22945 395
rect 5480 140 22945 150
rect 5480 120 5490 140
rect 5510 130 22945 140
rect 5510 120 5520 130
rect 5480 110 5520 120
rect 25415 105 25435 395
rect 28060 380 28100 390
rect 28060 370 28070 380
rect 5550 95 25435 105
rect 5550 75 5560 95
rect 5580 85 25435 95
rect 25460 360 28070 370
rect 28090 360 28100 380
rect 25460 350 28100 360
rect 5580 75 5590 85
rect 5550 65 5590 75
rect 1125 55 1165 65
rect 1125 35 1135 55
rect 1155 45 1165 55
rect 25460 45 25485 350
rect 30575 330 30595 395
rect 1155 35 25485 45
rect 1125 25 25485 35
rect 25505 310 30595 330
rect 1165 -10 1205 0
rect 1165 -30 1175 -10
rect 1195 -20 1205 -10
rect 25505 -20 25525 310
rect 33065 285 33090 395
rect 1195 -30 25525 -20
rect 1165 -40 25525 -30
rect 25545 265 33090 285
rect 25545 -60 25565 265
rect 35555 240 35575 395
rect 1275 -70 25565 -60
rect 1275 -90 1285 -70
rect 1305 -80 25565 -70
rect 25585 220 35575 240
rect 1305 -90 1315 -80
rect 1275 -100 1315 -90
rect 25585 -105 25605 220
rect 38045 195 38065 395
rect 1345 -115 25605 -105
rect 1345 -135 1355 -115
rect 1375 -125 25605 -115
rect 25625 175 38065 195
rect 1375 -135 1385 -125
rect 1345 -145 1385 -135
rect 25625 -150 25645 175
rect 40535 150 40555 395
rect 1410 -160 25645 -150
rect 1410 -180 1420 -160
rect 1440 -170 25645 -160
rect 25665 130 40555 150
rect 1440 -180 1450 -170
rect 1410 -190 1450 -180
rect 25665 -195 25685 130
rect 43025 105 43045 395
rect 1475 -205 25685 -195
rect 1475 -225 1485 -205
rect 1505 -215 25685 -205
rect 25705 85 43045 105
rect 1505 -225 1515 -215
rect 1475 -235 1515 -225
rect 25705 -240 25725 85
rect 45515 45 45535 395
rect 1545 -250 25725 -240
rect 1545 -270 1555 -250
rect 1575 -260 25725 -250
rect 25745 25 45535 45
rect 1575 -270 1585 -260
rect 1545 -280 1585 -270
rect 25745 -290 25765 25
rect 1615 -300 25765 -290
rect 1615 -320 1625 -300
rect 1645 -310 25765 -300
rect 1645 -320 1655 -310
rect 1615 -330 1655 -320
rect 125 -340 165 -330
rect 125 -360 135 -340
rect 155 -350 165 -340
rect 1255 -340 1295 -330
rect 1255 -350 1265 -340
rect 155 -360 1265 -350
rect 1285 -350 1295 -340
rect 2935 -340 2975 -330
rect 2935 -350 2945 -340
rect 1285 -360 2945 -350
rect 2965 -350 2975 -340
rect 4065 -340 4105 -330
rect 4065 -350 4075 -340
rect 2965 -360 4075 -350
rect 4095 -350 4105 -340
rect 5170 -340 5210 -330
rect 5170 -350 5180 -340
rect 4095 -360 5180 -350
rect 5200 -350 5210 -340
rect 6825 -340 6865 -330
rect 6825 -350 6835 -340
rect 5200 -360 6835 -350
rect 6855 -360 6865 -340
rect 125 -370 6865 -360
rect 55 -410 6775 -390
rect 55 -555 75 -410
rect 1165 -550 1185 -410
rect 2865 -550 2885 -410
rect 3995 -550 4015 -410
rect 5125 -550 5145 -410
rect 6755 -550 6775 -410
rect 3975 -570 3985 -550
rect 1125 -645 1360 -625
rect 1710 -645 1720 -625
rect 2250 -635 3060 -625
rect 1125 -1155 1145 -645
rect 2250 -655 2260 -635
rect 2280 -645 3060 -635
rect 3935 -645 4145 -625
rect 5065 -645 5295 -625
rect 6185 -635 6915 -625
rect 2280 -655 2290 -645
rect 2250 -665 2290 -655
rect 2250 -1145 2270 -665
rect 3935 -1135 3955 -645
rect 5065 -1130 5085 -645
rect 6185 -655 6195 -635
rect 6215 -645 6915 -635
rect 6215 -655 6225 -645
rect 6185 -665 6225 -655
rect 3930 -1150 3955 -1135
rect 5060 -1155 5085 -1130
rect 6190 -1140 6210 -665
rect 7845 -1125 7885 -1115
rect 7845 -1145 7855 -1125
rect 7875 -1145 7885 -1125
rect 7845 -1155 7885 -1145
rect 2315 -1285 2355 -1275
rect 2315 -1295 2325 -1285
rect 1135 -1315 1280 -1295
rect 2270 -1305 2325 -1295
rect 2345 -1295 2355 -1285
rect 6250 -1285 6290 -1275
rect 6250 -1295 6260 -1285
rect 2345 -1305 2970 -1295
rect 2270 -1315 2970 -1305
rect 3950 -1315 4100 -1295
rect 5070 -1315 5215 -1295
rect 6210 -1305 6260 -1295
rect 6280 -1295 6290 -1285
rect 8040 -1285 8080 -1275
rect 8040 -1295 8050 -1285
rect 6280 -1305 6855 -1295
rect 6210 -1315 6855 -1305
rect 7845 -1305 8050 -1295
rect 8070 -1305 8080 -1285
rect 7845 -1315 8080 -1305
rect 29375 -1410 29405 -1385
rect 30505 -1850 30540 -1830
rect 30520 -2145 30540 -1850
rect 33010 -2145 33030 -1835
rect 35485 -1860 35520 -1840
rect 37975 -1860 38010 -1840
rect 40455 -1860 40500 -1840
rect 42955 -1860 42990 -1840
rect 45445 -1860 45480 -1840
rect 47935 -1860 47970 -1840
rect 35500 -2145 35520 -1860
rect 37990 -2145 38010 -1860
rect 40480 -2145 40500 -1860
rect 42970 -2145 42990 -1860
rect 45460 -2145 45480 -1860
rect 47950 -2145 47970 -1860
rect 30365 -2155 30540 -2145
rect 30365 -2175 30375 -2155
rect 30395 -2165 30540 -2155
rect 32855 -2155 33030 -2145
rect 30395 -2175 30405 -2165
rect 2375 -2185 2415 -2175
rect 2375 -2195 2385 -2185
rect 1140 -2215 1275 -2195
rect 2270 -2205 2385 -2195
rect 2405 -2195 2415 -2185
rect 6310 -2185 6350 -2175
rect 6310 -2195 6320 -2185
rect 2405 -2205 2975 -2195
rect 2270 -2215 2975 -2205
rect 3955 -2215 4105 -2195
rect 5075 -2215 5220 -2195
rect 6210 -2205 6320 -2195
rect 6340 -2195 6350 -2185
rect 8085 -2185 8125 -2175
rect 30365 -2185 30405 -2175
rect 32855 -2175 32865 -2155
rect 32885 -2165 33030 -2155
rect 35345 -2155 35520 -2145
rect 32885 -2175 32895 -2165
rect 32855 -2185 32895 -2175
rect 35345 -2175 35355 -2155
rect 35375 -2165 35520 -2155
rect 37835 -2155 38010 -2145
rect 35375 -2175 35385 -2165
rect 35345 -2185 35385 -2175
rect 37835 -2175 37845 -2155
rect 37865 -2165 38010 -2155
rect 40325 -2155 40500 -2145
rect 37865 -2175 37875 -2165
rect 37835 -2185 37875 -2175
rect 40325 -2175 40335 -2155
rect 40355 -2165 40500 -2155
rect 42815 -2155 42990 -2145
rect 40355 -2175 40365 -2165
rect 40325 -2185 40365 -2175
rect 42815 -2175 42825 -2155
rect 42845 -2165 42990 -2155
rect 45305 -2155 45480 -2145
rect 42845 -2175 42855 -2165
rect 42815 -2185 42855 -2175
rect 45305 -2175 45315 -2155
rect 45335 -2165 45480 -2155
rect 47795 -2155 47970 -2145
rect 45335 -2175 45345 -2165
rect 45305 -2185 45345 -2175
rect 47795 -2175 47805 -2155
rect 47825 -2165 47970 -2155
rect 47825 -2175 47835 -2165
rect 47795 -2185 47835 -2175
rect 8085 -2195 8095 -2185
rect 6340 -2205 6855 -2195
rect 6210 -2215 6855 -2205
rect 7845 -2205 8095 -2195
rect 8115 -2205 8125 -2185
rect 7845 -2215 8125 -2205
rect 30550 -3075 30590 -3065
rect 2445 -3085 2485 -3075
rect 2445 -3095 2455 -3085
rect 1140 -3115 1275 -3095
rect 2270 -3105 2455 -3095
rect 2475 -3095 2485 -3085
rect 6380 -3085 6420 -3075
rect 6380 -3095 6390 -3085
rect 2475 -3105 2970 -3095
rect 2270 -3115 2970 -3105
rect 3950 -3115 4100 -3095
rect 5075 -3115 5220 -3095
rect 6210 -3105 6390 -3095
rect 6410 -3095 6420 -3085
rect 8135 -3085 8175 -3075
rect 8135 -3095 8145 -3085
rect 6410 -3105 6860 -3095
rect 6210 -3115 6860 -3105
rect 7845 -3105 8145 -3095
rect 8165 -3105 8175 -3085
rect 30550 -3095 30560 -3075
rect 30580 -3085 30590 -3075
rect 33040 -3075 33080 -3065
rect 30580 -3095 32940 -3085
rect 30550 -3105 32940 -3095
rect 33040 -3095 33050 -3075
rect 33070 -3085 33080 -3075
rect 35530 -3075 35570 -3065
rect 33070 -3095 35430 -3085
rect 33040 -3105 35430 -3095
rect 35530 -3095 35540 -3075
rect 35560 -3085 35570 -3075
rect 38020 -3075 38060 -3065
rect 35560 -3095 37920 -3085
rect 35530 -3105 37920 -3095
rect 38020 -3095 38030 -3075
rect 38050 -3085 38060 -3075
rect 40510 -3075 40550 -3065
rect 38050 -3095 40410 -3085
rect 38020 -3105 40410 -3095
rect 40510 -3095 40520 -3075
rect 40540 -3085 40550 -3075
rect 43000 -3075 43040 -3065
rect 40540 -3095 42900 -3085
rect 40510 -3105 42900 -3095
rect 43000 -3095 43010 -3075
rect 43030 -3080 43040 -3075
rect 45490 -3075 45530 -3065
rect 43030 -3085 43045 -3080
rect 43030 -3095 45390 -3085
rect 43000 -3105 45390 -3095
rect 45490 -3095 45500 -3075
rect 45520 -3085 45530 -3075
rect 45520 -3095 47880 -3085
rect 45490 -3105 47880 -3095
rect 7845 -3115 8175 -3105
rect 28060 -3120 28100 -3110
rect 28060 -3140 28070 -3120
rect 28090 -3130 28100 -3120
rect 28090 -3140 30455 -3130
rect 28060 -3150 30455 -3140
rect 30430 -3705 30455 -3150
rect 2510 -3985 2550 -3975
rect 2510 -3995 2520 -3985
rect 1140 -4015 1280 -3995
rect 1710 -4015 1830 -3995
rect 2270 -4005 2520 -3995
rect 2540 -3995 2550 -3985
rect 6445 -3985 6485 -3975
rect 6445 -3995 6455 -3985
rect 2540 -4005 2975 -3995
rect 2270 -4015 2975 -4005
rect 3950 -4015 4100 -3995
rect 5080 -4015 5225 -3995
rect 6210 -4005 6455 -3995
rect 6475 -3995 6485 -3985
rect 8185 -3985 8225 -3975
rect 8185 -3995 8195 -3985
rect 6475 -4005 6855 -3995
rect 6210 -4015 6855 -4005
rect 7845 -4005 8195 -3995
rect 8215 -4005 8225 -3985
rect 7845 -4015 8225 -4005
rect 25915 -4020 25955 -4010
rect 25915 -4025 25925 -4020
rect 25445 -4040 25925 -4025
rect 25945 -4040 25955 -4020
rect 25445 -4050 25955 -4040
rect 25445 -4435 25470 -4050
rect 25980 -4070 26020 -4060
rect 25980 -4075 25990 -4070
rect 10365 -4460 25470 -4435
rect 25495 -4090 25990 -4075
rect 26010 -4090 26020 -4070
rect 25495 -4100 26020 -4090
rect 8375 -4505 8415 -4495
rect 8375 -4525 8385 -4505
rect 8405 -4525 8415 -4505
rect 8375 -4535 8415 -4525
rect 8310 -4545 8350 -4535
rect 8310 -4565 8320 -4545
rect 8340 -4565 8350 -4545
rect 8310 -4575 8350 -4565
rect 8245 -4585 8285 -4575
rect 8245 -4595 8255 -4585
rect 7845 -4605 8255 -4595
rect 8275 -4605 8285 -4585
rect 7845 -4615 8285 -4605
rect 2575 -4885 2615 -4875
rect 2575 -4895 2585 -4885
rect 1130 -4915 1280 -4895
rect 1710 -4915 1835 -4895
rect 2270 -4905 2585 -4895
rect 2605 -4895 2615 -4885
rect 6510 -4885 6550 -4875
rect 6510 -4895 6520 -4885
rect 2605 -4905 2975 -4895
rect 2270 -4915 2975 -4905
rect 3940 -4915 4090 -4895
rect 5075 -4915 5220 -4895
rect 6210 -4905 6520 -4895
rect 6540 -4895 6550 -4885
rect 6540 -4905 6850 -4895
rect 6210 -4915 6850 -4905
rect 7845 -4915 7865 -4615
rect 8310 -4640 8330 -4575
rect 7890 -4660 8330 -4640
rect 2645 -5785 2685 -5775
rect 2645 -5795 2655 -5785
rect 1135 -5815 1275 -5795
rect 1710 -5815 1830 -5795
rect 2270 -5805 2655 -5795
rect 2675 -5795 2685 -5785
rect 6580 -5785 6620 -5775
rect 6580 -5795 6590 -5785
rect 2675 -5805 2965 -5795
rect 2270 -5815 2965 -5805
rect 3950 -5815 4100 -5795
rect 5080 -5815 5225 -5795
rect 6210 -5805 6590 -5795
rect 6610 -5795 6620 -5785
rect 7890 -5795 7910 -4660
rect 8375 -4685 8395 -4535
rect 6610 -5805 6855 -5795
rect 6210 -5815 6855 -5805
rect 7835 -5815 7910 -5795
rect 7935 -4705 8395 -4685
rect 7935 -6105 7955 -4705
rect 9245 -5025 9250 -5020
rect 10365 -5025 10385 -4460
rect 25495 -4485 25520 -4100
rect 26050 -4115 26090 -4105
rect 26050 -4120 26060 -4115
rect 12855 -4510 25520 -4485
rect 25540 -4135 26060 -4120
rect 26080 -4135 26090 -4115
rect 25540 -4145 26090 -4135
rect 12855 -5025 12875 -4510
rect 25540 -4535 25565 -4145
rect 26130 -4165 26170 -4155
rect 26130 -4170 26140 -4165
rect 15345 -4560 25565 -4535
rect 25585 -4185 26140 -4170
rect 26160 -4185 26170 -4165
rect 25585 -4195 26170 -4185
rect 15345 -5025 15365 -4560
rect 25585 -4585 25610 -4195
rect 26195 -4215 26235 -4205
rect 26195 -4220 26205 -4215
rect 17835 -4610 25610 -4585
rect 25630 -4235 26205 -4220
rect 26225 -4235 26235 -4215
rect 25630 -4245 26235 -4235
rect 17835 -5025 17855 -4610
rect 25630 -4640 25655 -4245
rect 26265 -4260 26305 -4250
rect 26265 -4265 26275 -4260
rect 20325 -4665 25655 -4640
rect 25680 -4280 26275 -4265
rect 26295 -4280 26305 -4260
rect 25680 -4290 26305 -4280
rect 25680 -4310 25710 -4290
rect 26335 -4305 26375 -4295
rect 26335 -4310 26345 -4305
rect 20325 -5025 20345 -4665
rect 25680 -4690 25705 -4310
rect 22815 -4715 25705 -4690
rect 25730 -4325 26345 -4310
rect 26365 -4325 26375 -4305
rect 25730 -4335 26375 -4325
rect 22815 -5025 22835 -4715
rect 25730 -4740 25755 -4335
rect 25305 -4765 25755 -4740
rect 27860 -4505 27900 -4495
rect 27860 -4525 27870 -4505
rect 27890 -4525 27900 -4505
rect 27860 -4535 27900 -4525
rect 25305 -5025 25325 -4765
rect 9310 -5045 9330 -5025
rect 10365 -5045 10450 -5025
rect 12855 -5045 12940 -5025
rect 15345 -5045 15430 -5025
rect 17835 -5045 17920 -5025
rect 20325 -5045 20410 -5025
rect 22815 -5045 22900 -5025
rect 25305 -5045 25390 -5025
rect 9305 -5050 9330 -5045
rect 9305 -5055 9325 -5050
rect 9300 -5220 9305 -5215
rect 9295 -5240 9305 -5220
rect 10430 -5485 10450 -5045
rect 12920 -5490 12940 -5045
rect 15410 -5495 15430 -5045
rect 17900 -5495 17920 -5045
rect 20390 -5495 20410 -5045
rect 22880 -5495 22900 -5045
rect 25370 -5495 25390 -5045
rect 27860 -5495 27885 -4535
rect 29375 -5040 29405 -5015
rect 30430 -5125 30450 -3705
rect 32920 -5125 32940 -3105
rect 35410 -5125 35430 -3105
rect 37900 -5125 37920 -3105
rect 40390 -5125 40410 -3105
rect 42880 -5125 42900 -3105
rect 45370 -5125 45390 -3105
rect 47860 -5125 47880 -3105
rect 30430 -5145 30540 -5125
rect 32920 -5145 33030 -5125
rect 35410 -5145 35520 -5125
rect 37900 -5145 38010 -5125
rect 40390 -5145 40500 -5125
rect 42880 -5145 42990 -5125
rect 45370 -5145 45480 -5125
rect 47860 -5145 47970 -5125
rect 30520 -5460 30540 -5145
rect 30505 -5480 30540 -5460
rect 33010 -5485 33030 -5145
rect 35500 -5470 35520 -5145
rect 37990 -5470 38010 -5145
rect 40480 -5470 40500 -5145
rect 42970 -5470 42990 -5145
rect 45460 -5470 45480 -5145
rect 47950 -5470 47970 -5145
rect 35485 -5490 35520 -5470
rect 37975 -5490 38010 -5470
rect 40465 -5490 40500 -5470
rect 42955 -5490 42990 -5470
rect 45445 -5490 45480 -5470
rect 47935 -5490 47970 -5470
rect 1120 -6535 1145 -6110
rect 2270 -6125 2780 -6105
rect 3930 -6125 3955 -6110
rect 2760 -6515 2780 -6125
rect 2740 -6525 2780 -6515
rect 1120 -6555 1380 -6535
rect 1710 -6555 1755 -6535
rect 2740 -6545 2750 -6525
rect 2770 -6535 2780 -6525
rect 3935 -6535 3955 -6125
rect 5065 -6535 5085 -6115
rect 6210 -6125 6715 -6105
rect 7835 -6125 7955 -6105
rect 6695 -6535 6715 -6125
rect 2770 -6545 3020 -6535
rect 2740 -6555 3020 -6545
rect 3935 -6555 4165 -6535
rect 5065 -6550 5305 -6535
rect 6675 -6545 6920 -6535
rect 5065 -6555 5280 -6550
rect 6675 -6565 6685 -6545
rect 6705 -6555 6920 -6545
rect 6705 -6565 6715 -6555
rect 6675 -6575 6715 -6565
rect 6185 -6685 6225 -6675
rect 6185 -6705 6195 -6685
rect 6215 -6695 6225 -6685
rect 6215 -6705 8025 -6695
rect 6185 -6715 7995 -6705
rect 7985 -6725 7995 -6715
rect 8015 -6715 8025 -6705
rect 10475 -6705 10515 -6695
rect 8015 -6725 8030 -6715
rect 7985 -6735 8030 -6725
rect 10475 -6725 10485 -6705
rect 10505 -6725 10515 -6705
rect 10475 -6735 10515 -6725
rect 12965 -6705 13005 -6695
rect 12965 -6725 12975 -6705
rect 12995 -6725 13005 -6705
rect 12965 -6735 13005 -6725
rect 15455 -6705 15495 -6695
rect 15455 -6725 15465 -6705
rect 15485 -6725 15495 -6705
rect 15455 -6735 15495 -6725
rect 17945 -6705 17985 -6695
rect 17945 -6725 17955 -6705
rect 17975 -6725 17985 -6705
rect 17945 -6735 17985 -6725
rect 20435 -6705 20475 -6695
rect 20435 -6725 20445 -6705
rect 20465 -6725 20475 -6705
rect 20435 -6735 20475 -6725
rect 22925 -6705 22965 -6695
rect 22925 -6725 22935 -6705
rect 22955 -6725 22965 -6705
rect 22925 -6735 22965 -6725
rect 25415 -6705 25455 -6695
rect 25415 -6725 25425 -6705
rect 25445 -6725 25455 -6705
rect 25415 -6735 25455 -6725
rect 30550 -6705 30590 -6695
rect 30550 -6725 30560 -6705
rect 30580 -6715 30590 -6705
rect 33040 -6705 33080 -6695
rect 30580 -6725 30595 -6715
rect 30550 -6735 30595 -6725
rect 33040 -6725 33050 -6705
rect 33070 -6710 33080 -6705
rect 35530 -6705 35570 -6695
rect 33070 -6725 33090 -6710
rect 33040 -6735 33090 -6725
rect 35530 -6725 35540 -6705
rect 35560 -6715 35570 -6705
rect 38020 -6705 38060 -6695
rect 35560 -6725 35575 -6715
rect 35530 -6735 35575 -6725
rect 38020 -6725 38030 -6705
rect 38050 -6715 38060 -6705
rect 40510 -6705 40550 -6695
rect 38050 -6725 38065 -6715
rect 38020 -6735 38065 -6725
rect 40510 -6725 40520 -6705
rect 40540 -6715 40550 -6705
rect 43000 -6705 43040 -6695
rect 40540 -6725 40555 -6715
rect 40510 -6735 40555 -6725
rect 43000 -6725 43010 -6705
rect 43030 -6710 43040 -6705
rect 45490 -6705 45530 -6695
rect 43030 -6725 43045 -6710
rect 43000 -6735 43045 -6725
rect 45490 -6725 45500 -6705
rect 45520 -6715 45530 -6705
rect 45520 -6725 45535 -6715
rect 45490 -6735 45535 -6725
rect 6225 -6750 6265 -6740
rect 6225 -6770 6235 -6750
rect 6255 -6760 6265 -6750
rect 10475 -6760 10495 -6735
rect 6255 -6770 10495 -6760
rect 6225 -6780 10495 -6770
rect 12965 -6800 12990 -6735
rect 6335 -6810 12990 -6800
rect 6335 -6830 6345 -6810
rect 6365 -6820 12990 -6810
rect 6365 -6830 6375 -6820
rect 6335 -6840 6375 -6830
rect 15455 -6845 15475 -6735
rect 6405 -6855 15475 -6845
rect 6405 -6875 6415 -6855
rect 6435 -6865 15475 -6855
rect 6435 -6875 6445 -6865
rect 6405 -6885 6445 -6875
rect 17945 -6890 17965 -6735
rect 6470 -6900 17965 -6890
rect 6470 -6920 6480 -6900
rect 6500 -6910 17965 -6900
rect 6500 -6920 6510 -6910
rect 6470 -6930 6510 -6920
rect 20435 -6935 20455 -6735
rect 6535 -6945 20455 -6935
rect 6535 -6965 6545 -6945
rect 6565 -6955 20455 -6945
rect 6565 -6965 6575 -6955
rect 6535 -6975 6575 -6965
rect 22925 -6980 22945 -6735
rect 6605 -6990 22945 -6980
rect 6605 -7010 6615 -6990
rect 6635 -7000 22945 -6990
rect 6635 -7010 6645 -7000
rect 6605 -7020 6645 -7010
rect 25415 -7025 25435 -6735
rect 28060 -6750 28100 -6740
rect 28060 -6760 28070 -6750
rect 6675 -7035 25435 -7025
rect 6675 -7055 6685 -7035
rect 6705 -7045 25435 -7035
rect 25460 -6770 28070 -6760
rect 28090 -6770 28100 -6750
rect 25460 -6780 28100 -6770
rect 6705 -7055 6715 -7045
rect 6675 -7065 6715 -7055
rect 2250 -7075 2290 -7065
rect 2250 -7095 2260 -7075
rect 2280 -7085 2290 -7075
rect 25460 -7085 25485 -6780
rect 30575 -6800 30595 -6735
rect 2280 -7095 25485 -7085
rect 2250 -7105 25485 -7095
rect 25505 -6820 30595 -6800
rect 2290 -7140 2330 -7130
rect 2290 -7160 2300 -7140
rect 2320 -7150 2330 -7140
rect 25505 -7150 25525 -6820
rect 33065 -6845 33090 -6735
rect 2320 -7160 25525 -7150
rect 2290 -7170 25525 -7160
rect 25545 -6865 33090 -6845
rect 25545 -7190 25565 -6865
rect 35555 -6890 35575 -6735
rect 2400 -7200 25565 -7190
rect 2400 -7220 2410 -7200
rect 2430 -7210 25565 -7200
rect 25585 -6910 35575 -6890
rect 2430 -7220 2440 -7210
rect 2400 -7230 2440 -7220
rect 25585 -7235 25605 -6910
rect 38045 -6935 38065 -6735
rect 2470 -7245 25605 -7235
rect 2470 -7265 2480 -7245
rect 2500 -7255 25605 -7245
rect 25625 -6955 38065 -6935
rect 2500 -7265 2510 -7255
rect 2470 -7275 2510 -7265
rect 25625 -7280 25645 -6955
rect 40535 -6980 40555 -6735
rect 2535 -7290 25645 -7280
rect 2535 -7310 2545 -7290
rect 2565 -7300 25645 -7290
rect 25665 -7000 40555 -6980
rect 2565 -7310 2575 -7300
rect 2535 -7320 2575 -7310
rect 25665 -7325 25685 -7000
rect 43025 -7025 43045 -6735
rect 2600 -7335 25685 -7325
rect 2600 -7355 2610 -7335
rect 2630 -7345 25685 -7335
rect 25705 -7045 43045 -7025
rect 2630 -7355 2640 -7345
rect 2600 -7365 2640 -7355
rect 25705 -7370 25725 -7045
rect 45515 -7085 45535 -6735
rect 2670 -7380 25725 -7370
rect 2670 -7400 2680 -7380
rect 2700 -7390 25725 -7380
rect 25745 -7105 45535 -7085
rect 2700 -7400 2710 -7390
rect 2670 -7410 2710 -7400
rect 25745 -7420 25765 -7105
rect 2740 -7430 25765 -7420
rect 2740 -7450 2750 -7430
rect 2770 -7440 25765 -7430
rect 2770 -7450 2780 -7440
rect 2740 -7460 2780 -7450
rect 125 -7480 165 -7470
rect 125 -7500 135 -7480
rect 155 -7490 165 -7480
rect 1255 -7480 1295 -7470
rect 1255 -7490 1265 -7480
rect 155 -7500 1265 -7490
rect 1285 -7490 1295 -7480
rect 2935 -7480 2975 -7470
rect 2935 -7490 2945 -7480
rect 1285 -7500 2945 -7490
rect 2965 -7490 2975 -7480
rect 4065 -7480 4105 -7470
rect 4065 -7490 4075 -7480
rect 2965 -7500 4075 -7490
rect 4095 -7490 4105 -7480
rect 5170 -7480 5210 -7470
rect 5170 -7490 5180 -7480
rect 4095 -7500 5180 -7490
rect 5200 -7490 5210 -7480
rect 6825 -7480 6865 -7470
rect 6825 -7490 6835 -7480
rect 5200 -7500 6835 -7490
rect 6855 -7500 6865 -7480
rect 125 -7510 6865 -7500
rect 55 -7550 6775 -7530
rect 55 -7695 75 -7550
rect 1165 -7690 1185 -7550
rect 2865 -7690 2885 -7550
rect 3995 -7690 4015 -7550
rect 5125 -7690 5145 -7550
rect 6755 -7690 6775 -7550
rect 3975 -7710 3985 -7690
rect 1125 -7785 1360 -7765
rect 1710 -7785 1720 -7765
rect 2250 -7775 3060 -7765
rect 1125 -8295 1145 -7785
rect 2250 -7795 2260 -7775
rect 2280 -7785 3060 -7775
rect 3935 -7785 4145 -7765
rect 5065 -7785 5295 -7765
rect 6185 -7775 6915 -7765
rect 2280 -7795 2290 -7785
rect 2250 -7805 2290 -7795
rect 2250 -8285 2270 -7805
rect 3935 -8275 3955 -7785
rect 5065 -8270 5085 -7785
rect 6185 -7795 6195 -7775
rect 6215 -7785 6915 -7775
rect 6215 -7795 6225 -7785
rect 6185 -7805 6225 -7795
rect 3930 -8290 3955 -8275
rect 5060 -8295 5085 -8270
rect 6190 -8280 6210 -7805
rect 30355 -8155 30415 -8135
rect 30355 -8175 30375 -8155
rect 30395 -8175 30415 -8155
rect 30355 -8195 30415 -8175
rect 32845 -8155 32905 -8135
rect 32845 -8175 32865 -8155
rect 32885 -8175 32905 -8155
rect 32845 -8195 32905 -8175
rect 35335 -8155 35395 -8135
rect 35335 -8175 35355 -8155
rect 35375 -8175 35395 -8155
rect 35335 -8195 35395 -8175
rect 37825 -8155 37885 -8135
rect 37825 -8175 37845 -8155
rect 37865 -8175 37885 -8155
rect 37825 -8195 37885 -8175
rect 40315 -8155 40375 -8135
rect 40315 -8175 40335 -8155
rect 40355 -8175 40375 -8155
rect 40315 -8195 40375 -8175
rect 42805 -8155 42865 -8135
rect 42805 -8175 42825 -8155
rect 42845 -8175 42865 -8155
rect 42805 -8195 42865 -8175
rect 45295 -8155 45355 -8135
rect 45295 -8175 45315 -8155
rect 45335 -8175 45355 -8155
rect 45295 -8195 45355 -8175
rect 47785 -8155 47845 -8135
rect 47785 -8175 47805 -8155
rect 47825 -8175 47845 -8155
rect 47785 -8195 47845 -8175
rect 30355 -8215 30375 -8195
rect 32845 -8215 32865 -8195
rect 35335 -8215 35355 -8195
rect 37825 -8215 37845 -8195
rect 40315 -8215 40335 -8195
rect 42805 -8215 42825 -8195
rect 45295 -8215 45315 -8195
rect 47785 -8215 47805 -8195
rect 30345 -8225 30385 -8215
rect 30345 -8245 30355 -8225
rect 30375 -8245 30385 -8225
rect 30345 -8255 30385 -8245
rect 32835 -8225 32875 -8215
rect 32835 -8245 32845 -8225
rect 32865 -8245 32875 -8225
rect 32835 -8255 32875 -8245
rect 35325 -8225 35365 -8215
rect 35325 -8245 35335 -8225
rect 35355 -8245 35365 -8225
rect 35325 -8255 35365 -8245
rect 37815 -8225 37855 -8215
rect 37815 -8245 37825 -8225
rect 37845 -8245 37855 -8225
rect 37815 -8255 37855 -8245
rect 40305 -8225 40345 -8215
rect 40305 -8245 40315 -8225
rect 40335 -8245 40345 -8225
rect 40305 -8255 40345 -8245
rect 42795 -8225 42835 -8215
rect 42795 -8245 42805 -8225
rect 42825 -8245 42835 -8225
rect 42795 -8255 42835 -8245
rect 45285 -8225 45325 -8215
rect 45285 -8245 45295 -8225
rect 45315 -8245 45325 -8225
rect 45285 -8255 45325 -8245
rect 47775 -8225 47815 -8215
rect 47775 -8245 47785 -8225
rect 47805 -8245 47815 -8225
rect 47775 -8255 47815 -8245
rect 7845 -8265 7885 -8255
rect 7845 -8285 7855 -8265
rect 7875 -8285 7885 -8265
rect 7845 -8295 7885 -8285
rect 2315 -8425 2355 -8415
rect 2315 -8435 2325 -8425
rect 1135 -8455 1280 -8435
rect 2270 -8445 2325 -8435
rect 2345 -8435 2355 -8425
rect 6250 -8425 6290 -8415
rect 6250 -8435 6260 -8425
rect 2345 -8445 2970 -8435
rect 2270 -8455 2970 -8445
rect 3950 -8455 4100 -8435
rect 5070 -8455 5215 -8435
rect 6210 -8445 6260 -8435
rect 6280 -8435 6290 -8425
rect 8040 -8425 8080 -8415
rect 8040 -8435 8050 -8425
rect 6280 -8445 6855 -8435
rect 6210 -8455 6855 -8445
rect 7845 -8445 8050 -8435
rect 8070 -8445 8080 -8425
rect 7845 -8455 8080 -8445
rect 29375 -8930 29405 -8905
rect 2375 -9325 2415 -9315
rect 2375 -9335 2385 -9325
rect 1140 -9355 1275 -9335
rect 2270 -9345 2385 -9335
rect 2405 -9335 2415 -9325
rect 6310 -9325 6350 -9315
rect 6310 -9335 6320 -9325
rect 2405 -9345 2975 -9335
rect 2270 -9355 2975 -9345
rect 3955 -9355 4105 -9335
rect 5075 -9355 5220 -9335
rect 6210 -9345 6320 -9335
rect 6340 -9335 6350 -9325
rect 8085 -9325 8125 -9315
rect 8085 -9335 8095 -9325
rect 6340 -9345 6855 -9335
rect 6210 -9355 6855 -9345
rect 7845 -9345 8095 -9335
rect 8115 -9345 8125 -9325
rect 7845 -9355 8125 -9345
rect 2445 -10225 2485 -10215
rect 2445 -10235 2455 -10225
rect 1140 -10255 1275 -10235
rect 2270 -10245 2455 -10235
rect 2475 -10235 2485 -10225
rect 6380 -10225 6420 -10215
rect 6380 -10235 6390 -10225
rect 2475 -10245 2970 -10235
rect 2270 -10255 2970 -10245
rect 3950 -10255 4100 -10235
rect 5075 -10255 5220 -10235
rect 6210 -10245 6390 -10235
rect 6410 -10235 6420 -10225
rect 8135 -10225 8175 -10215
rect 8135 -10235 8145 -10225
rect 6410 -10245 6860 -10235
rect 6210 -10255 6860 -10245
rect 7845 -10245 8145 -10235
rect 8165 -10245 8175 -10225
rect 7845 -10255 8175 -10245
rect 30550 -10595 30590 -10585
rect 30550 -10615 30560 -10595
rect 30580 -10605 30590 -10595
rect 33040 -10595 33080 -10585
rect 30580 -10615 32945 -10605
rect 30550 -10625 32945 -10615
rect 33040 -10615 33050 -10595
rect 33070 -10600 33080 -10595
rect 35530 -10595 35570 -10585
rect 33070 -10605 33090 -10600
rect 33070 -10615 35435 -10605
rect 33040 -10625 35435 -10615
rect 35530 -10615 35540 -10595
rect 35560 -10605 35570 -10595
rect 38020 -10595 38060 -10585
rect 35560 -10615 37925 -10605
rect 35530 -10625 37925 -10615
rect 38020 -10615 38030 -10595
rect 38050 -10605 38060 -10595
rect 40510 -10595 40550 -10585
rect 38050 -10615 40415 -10605
rect 38020 -10625 40415 -10615
rect 40510 -10615 40520 -10595
rect 40540 -10605 40550 -10595
rect 43000 -10595 43040 -10585
rect 40540 -10615 42905 -10605
rect 40510 -10625 42905 -10615
rect 43000 -10615 43010 -10595
rect 43030 -10600 43040 -10595
rect 45490 -10595 45530 -10585
rect 43030 -10605 43045 -10600
rect 43030 -10615 45395 -10605
rect 43000 -10625 45395 -10615
rect 45490 -10615 45500 -10595
rect 45520 -10605 45530 -10595
rect 45520 -10615 47885 -10605
rect 45490 -10625 47885 -10615
rect 28060 -10640 28100 -10630
rect 28060 -10660 28070 -10640
rect 28090 -10650 28100 -10640
rect 28090 -10660 30455 -10650
rect 28060 -10670 30455 -10660
rect 2510 -11125 2550 -11115
rect 2510 -11135 2520 -11125
rect 1140 -11155 1280 -11135
rect 1710 -11155 1830 -11135
rect 2270 -11145 2520 -11135
rect 2540 -11135 2550 -11125
rect 6445 -11125 6485 -11115
rect 6445 -11135 6455 -11125
rect 2540 -11145 2975 -11135
rect 2270 -11155 2975 -11145
rect 3950 -11155 4100 -11135
rect 5080 -11155 5225 -11135
rect 6210 -11145 6455 -11135
rect 6475 -11135 6485 -11125
rect 8185 -11125 8225 -11115
rect 8185 -11135 8195 -11125
rect 6475 -11145 6855 -11135
rect 6210 -11155 6855 -11145
rect 7845 -11145 8195 -11135
rect 8215 -11145 8225 -11125
rect 7845 -11155 8225 -11145
rect 25915 -11160 25955 -11150
rect 25915 -11165 25925 -11160
rect 25445 -11180 25925 -11165
rect 25945 -11180 25955 -11160
rect 25445 -11190 25955 -11180
rect 25445 -11575 25470 -11190
rect 25980 -11210 26020 -11200
rect 25980 -11215 25990 -11210
rect 10365 -11600 25470 -11575
rect 25495 -11230 25990 -11215
rect 26010 -11230 26020 -11210
rect 25495 -11240 26020 -11230
rect 8375 -11645 8415 -11635
rect 8375 -11665 8385 -11645
rect 8405 -11665 8415 -11645
rect 8375 -11675 8415 -11665
rect 8310 -11685 8350 -11675
rect 8310 -11705 8320 -11685
rect 8340 -11705 8350 -11685
rect 8310 -11715 8350 -11705
rect 8245 -11725 8285 -11715
rect 8245 -11735 8255 -11725
rect 7845 -11745 8255 -11735
rect 8275 -11745 8285 -11725
rect 7845 -11755 8285 -11745
rect 2575 -12025 2615 -12015
rect 2575 -12035 2585 -12025
rect 1130 -12055 1280 -12035
rect 1710 -12055 1835 -12035
rect 2270 -12045 2585 -12035
rect 2605 -12035 2615 -12025
rect 6510 -12025 6550 -12015
rect 6510 -12035 6520 -12025
rect 2605 -12045 2975 -12035
rect 2270 -12055 2975 -12045
rect 3940 -12055 4090 -12035
rect 5075 -12055 5220 -12035
rect 6210 -12045 6520 -12035
rect 6540 -12035 6550 -12025
rect 6540 -12045 6850 -12035
rect 6210 -12055 6850 -12045
rect 7845 -12055 7865 -11755
rect 8310 -11780 8330 -11715
rect 7890 -11800 8330 -11780
rect 2645 -12925 2685 -12915
rect 2645 -12935 2655 -12925
rect 1135 -12955 1275 -12935
rect 1710 -12955 1830 -12935
rect 2270 -12945 2655 -12935
rect 2675 -12935 2685 -12925
rect 6580 -12925 6620 -12915
rect 6580 -12935 6590 -12925
rect 2675 -12945 2965 -12935
rect 2270 -12955 2965 -12945
rect 3950 -12955 4100 -12935
rect 5080 -12955 5225 -12935
rect 6210 -12945 6590 -12935
rect 6610 -12935 6620 -12925
rect 7890 -12935 7910 -11800
rect 8375 -11825 8395 -11675
rect 6610 -12945 6855 -12935
rect 6210 -12955 6855 -12945
rect 7835 -12955 7910 -12935
rect 7935 -11845 8395 -11825
rect 7935 -13245 7955 -11845
rect 9245 -12165 9250 -12160
rect 10365 -12165 10385 -11600
rect 25495 -11625 25520 -11240
rect 26050 -11255 26090 -11245
rect 26050 -11260 26060 -11255
rect 12855 -11650 25520 -11625
rect 25540 -11275 26060 -11260
rect 26080 -11275 26090 -11255
rect 25540 -11285 26090 -11275
rect 12855 -12165 12875 -11650
rect 25540 -11675 25565 -11285
rect 26130 -11305 26170 -11295
rect 26130 -11310 26140 -11305
rect 15345 -11700 25565 -11675
rect 25585 -11325 26140 -11310
rect 26160 -11325 26170 -11305
rect 25585 -11335 26170 -11325
rect 15345 -12165 15365 -11700
rect 25585 -11725 25610 -11335
rect 26195 -11355 26235 -11345
rect 26195 -11360 26205 -11355
rect 17835 -11750 25610 -11725
rect 25630 -11375 26205 -11360
rect 26225 -11375 26235 -11355
rect 25630 -11385 26235 -11375
rect 17835 -12165 17855 -11750
rect 25630 -11780 25655 -11385
rect 26265 -11400 26305 -11390
rect 26265 -11405 26275 -11400
rect 20325 -11805 25655 -11780
rect 25680 -11420 26275 -11405
rect 26295 -11420 26305 -11400
rect 25680 -11430 26305 -11420
rect 25680 -11450 25710 -11430
rect 26335 -11445 26375 -11435
rect 26335 -11450 26345 -11445
rect 20325 -12165 20345 -11805
rect 25680 -11830 25705 -11450
rect 22815 -11855 25705 -11830
rect 25730 -11465 26345 -11450
rect 26365 -11465 26375 -11445
rect 25730 -11475 26375 -11465
rect 22815 -12165 22835 -11855
rect 25730 -11880 25755 -11475
rect 25305 -11905 25755 -11880
rect 27860 -11645 27900 -11635
rect 27860 -11665 27870 -11645
rect 27890 -11665 27900 -11645
rect 27860 -11675 27900 -11665
rect 25305 -12165 25325 -11905
rect 9310 -12185 9330 -12165
rect 10365 -12185 10450 -12165
rect 12855 -12185 12940 -12165
rect 15345 -12185 15430 -12165
rect 17835 -12185 17920 -12165
rect 20325 -12185 20410 -12165
rect 22815 -12185 22900 -12165
rect 25305 -12185 25390 -12165
rect 9305 -12190 9330 -12185
rect 9305 -12195 9325 -12190
rect 9300 -12360 9305 -12355
rect 9295 -12380 9305 -12360
rect 10430 -12625 10450 -12185
rect 12920 -12630 12940 -12185
rect 15410 -12635 15430 -12185
rect 17900 -12635 17920 -12185
rect 20390 -12635 20410 -12185
rect 22880 -12635 22900 -12185
rect 25370 -12635 25390 -12185
rect 27860 -12635 27885 -11675
rect 29375 -12180 29405 -12155
rect 30435 -12165 30455 -10670
rect 30435 -12185 30540 -12165
rect 30520 -12600 30540 -12185
rect 32925 -12175 32945 -10625
rect 35415 -12175 35435 -10625
rect 37905 -12175 37925 -10625
rect 40395 -12175 40415 -10625
rect 42885 -12175 42905 -10625
rect 45375 -12175 45395 -10625
rect 47865 -12175 47885 -10625
rect 32925 -12195 33030 -12175
rect 35415 -12195 35520 -12175
rect 37905 -12195 38010 -12175
rect 40395 -12195 40500 -12175
rect 42885 -12195 42990 -12175
rect 45375 -12195 45480 -12175
rect 47865 -12195 47970 -12175
rect 30500 -12620 30540 -12600
rect 33010 -12625 33030 -12195
rect 35500 -12610 35520 -12195
rect 37990 -12610 38010 -12195
rect 40480 -12610 40500 -12195
rect 42970 -12610 42990 -12195
rect 45460 -12610 45480 -12195
rect 47950 -12610 47970 -12195
rect 35485 -12630 35520 -12610
rect 37975 -12630 38010 -12610
rect 40460 -12630 40500 -12610
rect 42950 -12630 42990 -12610
rect 45440 -12630 45480 -12610
rect 47935 -12630 47970 -12610
rect 1120 -13675 1145 -13250
rect 2270 -13265 2780 -13245
rect 3930 -13265 3955 -13250
rect 2760 -13655 2780 -13265
rect 2740 -13665 2780 -13655
rect 1120 -13695 1380 -13675
rect 1710 -13695 1755 -13675
rect 2740 -13685 2750 -13665
rect 2770 -13675 2780 -13665
rect 3935 -13675 3955 -13265
rect 5065 -13675 5085 -13255
rect 6210 -13265 6715 -13245
rect 7835 -13265 7955 -13245
rect 6695 -13675 6715 -13265
rect 2770 -13685 3020 -13675
rect 2740 -13695 3020 -13685
rect 3935 -13695 4165 -13675
rect 5065 -13690 5305 -13675
rect 6675 -13685 6920 -13675
rect 5065 -13695 5280 -13690
rect 6675 -13705 6685 -13685
rect 6705 -13695 6920 -13685
rect 6705 -13705 6715 -13695
rect 6675 -13715 6715 -13705
rect 6185 -13825 6225 -13815
rect 6185 -13845 6195 -13825
rect 6215 -13835 6225 -13825
rect 6215 -13845 8025 -13835
rect 6185 -13855 7995 -13845
rect 7985 -13865 7995 -13855
rect 8015 -13855 8025 -13845
rect 10475 -13845 10515 -13835
rect 8015 -13865 8030 -13855
rect 7985 -13875 8030 -13865
rect 10475 -13865 10485 -13845
rect 10505 -13865 10515 -13845
rect 10475 -13875 10515 -13865
rect 12965 -13845 13005 -13835
rect 12965 -13865 12975 -13845
rect 12995 -13865 13005 -13845
rect 12965 -13875 13005 -13865
rect 15455 -13845 15495 -13835
rect 15455 -13865 15465 -13845
rect 15485 -13865 15495 -13845
rect 15455 -13875 15495 -13865
rect 17945 -13845 17985 -13835
rect 17945 -13865 17955 -13845
rect 17975 -13865 17985 -13845
rect 17945 -13875 17985 -13865
rect 20435 -13845 20475 -13835
rect 20435 -13865 20445 -13845
rect 20465 -13865 20475 -13845
rect 20435 -13875 20475 -13865
rect 22925 -13845 22965 -13835
rect 22925 -13865 22935 -13845
rect 22955 -13865 22965 -13845
rect 22925 -13875 22965 -13865
rect 25415 -13845 25455 -13835
rect 25415 -13865 25425 -13845
rect 25445 -13865 25455 -13845
rect 25415 -13875 25455 -13865
rect 30550 -13845 30590 -13835
rect 30550 -13865 30560 -13845
rect 30580 -13855 30590 -13845
rect 33040 -13845 33080 -13835
rect 30580 -13865 30595 -13855
rect 30550 -13875 30595 -13865
rect 33040 -13865 33050 -13845
rect 33070 -13850 33080 -13845
rect 35530 -13845 35570 -13835
rect 33070 -13865 33090 -13850
rect 33040 -13875 33090 -13865
rect 35530 -13865 35540 -13845
rect 35560 -13855 35570 -13845
rect 38020 -13845 38060 -13835
rect 35560 -13865 35575 -13855
rect 35530 -13875 35575 -13865
rect 38020 -13865 38030 -13845
rect 38050 -13855 38060 -13845
rect 40510 -13845 40550 -13835
rect 38050 -13865 38065 -13855
rect 38020 -13875 38065 -13865
rect 40510 -13865 40520 -13845
rect 40540 -13855 40550 -13845
rect 43000 -13845 43040 -13835
rect 40540 -13865 40555 -13855
rect 40510 -13875 40555 -13865
rect 43000 -13865 43010 -13845
rect 43030 -13850 43040 -13845
rect 45490 -13845 45530 -13835
rect 43030 -13865 43045 -13850
rect 43000 -13875 43045 -13865
rect 45490 -13865 45500 -13845
rect 45520 -13855 45530 -13845
rect 45520 -13865 45535 -13855
rect 45490 -13875 45535 -13865
rect 6225 -13890 6265 -13880
rect 6225 -13910 6235 -13890
rect 6255 -13900 6265 -13890
rect 10475 -13900 10495 -13875
rect 6255 -13910 10495 -13900
rect 6225 -13920 10495 -13910
rect 12965 -13940 12990 -13875
rect 6335 -13950 12990 -13940
rect 6335 -13970 6345 -13950
rect 6365 -13960 12990 -13950
rect 6365 -13970 6375 -13960
rect 6335 -13980 6375 -13970
rect 15455 -13985 15475 -13875
rect 6405 -13995 15475 -13985
rect 6405 -14015 6415 -13995
rect 6435 -14005 15475 -13995
rect 6435 -14015 6445 -14005
rect 6405 -14025 6445 -14015
rect 17945 -14030 17965 -13875
rect 6470 -14040 17965 -14030
rect 6470 -14060 6480 -14040
rect 6500 -14050 17965 -14040
rect 6500 -14060 6510 -14050
rect 6470 -14070 6510 -14060
rect 20435 -14075 20455 -13875
rect 6535 -14085 20455 -14075
rect 6535 -14105 6545 -14085
rect 6565 -14095 20455 -14085
rect 6565 -14105 6575 -14095
rect 6535 -14115 6575 -14105
rect 22925 -14120 22945 -13875
rect 6605 -14130 22945 -14120
rect 6605 -14150 6615 -14130
rect 6635 -14140 22945 -14130
rect 6635 -14150 6645 -14140
rect 6605 -14160 6645 -14150
rect 25415 -14165 25435 -13875
rect 28060 -13890 28100 -13880
rect 28060 -13900 28070 -13890
rect 6675 -14175 25435 -14165
rect 6675 -14195 6685 -14175
rect 6705 -14185 25435 -14175
rect 25460 -13910 28070 -13900
rect 28090 -13910 28100 -13890
rect 25460 -13920 28100 -13910
rect 6705 -14195 6715 -14185
rect 6675 -14205 6715 -14195
rect 2250 -14215 2290 -14205
rect 2250 -14235 2260 -14215
rect 2280 -14225 2290 -14215
rect 25460 -14225 25485 -13920
rect 30575 -13940 30595 -13875
rect 2280 -14235 25485 -14225
rect 2250 -14245 25485 -14235
rect 25505 -13960 30595 -13940
rect 2290 -14280 2330 -14270
rect 2290 -14300 2300 -14280
rect 2320 -14290 2330 -14280
rect 25505 -14290 25525 -13960
rect 33065 -13985 33090 -13875
rect 2320 -14300 25525 -14290
rect 2290 -14310 25525 -14300
rect 25545 -14005 33090 -13985
rect 25545 -14330 25565 -14005
rect 35555 -14030 35575 -13875
rect 2400 -14340 25565 -14330
rect 2400 -14360 2410 -14340
rect 2430 -14350 25565 -14340
rect 25585 -14050 35575 -14030
rect 2430 -14360 2440 -14350
rect 2400 -14370 2440 -14360
rect 25585 -14375 25605 -14050
rect 38045 -14075 38065 -13875
rect 2470 -14385 25605 -14375
rect 2470 -14405 2480 -14385
rect 2500 -14395 25605 -14385
rect 25625 -14095 38065 -14075
rect 2500 -14405 2510 -14395
rect 2470 -14415 2510 -14405
rect 25625 -14420 25645 -14095
rect 40535 -14120 40555 -13875
rect 2535 -14430 25645 -14420
rect 2535 -14450 2545 -14430
rect 2565 -14440 25645 -14430
rect 25665 -14140 40555 -14120
rect 2565 -14450 2575 -14440
rect 2535 -14460 2575 -14450
rect 25665 -14465 25685 -14140
rect 43025 -14165 43045 -13875
rect 2600 -14475 25685 -14465
rect 2600 -14495 2610 -14475
rect 2630 -14485 25685 -14475
rect 25705 -14185 43045 -14165
rect 2630 -14495 2640 -14485
rect 2600 -14505 2640 -14495
rect 25705 -14510 25725 -14185
rect 45515 -14225 45535 -13875
rect 2670 -14520 25725 -14510
rect 2670 -14540 2680 -14520
rect 2700 -14530 25725 -14520
rect 25745 -14245 45535 -14225
rect 2700 -14540 2710 -14530
rect 2670 -14550 2710 -14540
rect 25745 -14560 25765 -14245
rect 2740 -14570 25765 -14560
rect 2740 -14590 2750 -14570
rect 2770 -14580 25765 -14570
rect 2770 -14590 2780 -14580
rect 2740 -14600 2780 -14590
<< viali >>
rect 30375 -2175 30395 -2155
rect 32865 -2175 32885 -2155
rect 35355 -2175 35375 -2155
rect 37845 -2175 37865 -2155
rect 40335 -2175 40355 -2155
rect 42825 -2175 42845 -2155
rect 45315 -2175 45335 -2155
rect 47805 -2175 47825 -2155
rect 30375 -8175 30395 -8155
rect 32865 -8175 32885 -8155
rect 35355 -8175 35375 -8155
rect 37845 -8175 37865 -8155
rect 40335 -8175 40355 -8155
rect 42825 -8175 42845 -8155
rect 45315 -8175 45335 -8155
rect 47805 -8175 47825 -8155
<< metal1 >>
rect 605 6305 1895 6405
rect 2285 6305 3025 6405
rect 3415 6305 4455 6405
rect 4545 6305 6900 6405
rect 7825 1995 8105 2085
rect 7890 1685 8110 1775
rect 7890 1455 7995 1685
rect 27845 1675 28190 1780
rect 7830 1355 7995 1455
rect 27855 1380 28255 1480
rect 625 750 865 850
rect 730 -725 865 750
rect 27870 780 28180 885
rect 1730 -725 2055 -720
rect 605 -815 1725 -725
rect 1730 -815 3025 -725
rect 605 -825 3025 -815
rect 3415 -825 4455 -725
rect 4545 -825 5290 -725
rect 5670 -820 6900 -725
rect 5790 -825 6900 -820
rect 1075 -830 3010 -825
rect 27870 -1720 28005 780
rect 27870 -1830 28190 -1720
rect 27945 -2120 28255 -2020
rect 30355 -2145 30415 -2135
rect 30355 -2185 30365 -2145
rect 30405 -2185 30415 -2145
rect 30355 -2195 30415 -2185
rect 32845 -2145 32905 -2135
rect 32845 -2185 32855 -2145
rect 32895 -2185 32905 -2145
rect 32845 -2195 32905 -2185
rect 35335 -2145 35395 -2135
rect 35335 -2185 35345 -2145
rect 35385 -2185 35395 -2145
rect 35335 -2195 35395 -2185
rect 37825 -2145 37885 -2135
rect 37825 -2185 37835 -2145
rect 37875 -2185 37885 -2145
rect 37825 -2195 37885 -2185
rect 40315 -2145 40375 -2135
rect 40315 -2185 40325 -2145
rect 40365 -2185 40375 -2145
rect 40315 -2195 40375 -2185
rect 42805 -2145 42865 -2135
rect 42805 -2185 42815 -2145
rect 42855 -2185 42865 -2145
rect 42805 -2195 42865 -2185
rect 45295 -2145 45355 -2135
rect 45295 -2185 45305 -2145
rect 45345 -2185 45355 -2145
rect 45295 -2195 45355 -2185
rect 47785 -2145 47845 -2135
rect 47785 -2185 47795 -2145
rect 47835 -2185 47845 -2145
rect 47785 -2195 47845 -2185
rect 7825 -5135 8105 -5045
rect 7890 -5445 8110 -5355
rect 7890 -5675 7995 -5445
rect 27845 -5455 28190 -5350
rect 7830 -5775 7995 -5675
rect 27855 -5750 28255 -5650
rect 615 -6375 845 -6280
rect 730 -7470 845 -6375
rect 730 -7865 865 -7470
rect 1730 -7865 2055 -7860
rect 605 -7955 1725 -7865
rect 1730 -7955 3025 -7865
rect 605 -7965 3025 -7955
rect 3415 -7965 4455 -7865
rect 4545 -7965 5290 -7865
rect 5670 -7960 6900 -7865
rect 5790 -7965 6900 -7960
rect 1075 -7970 3010 -7965
rect 30355 -8145 30415 -8135
rect 30355 -8185 30365 -8145
rect 30405 -8185 30415 -8145
rect 30355 -8195 30415 -8185
rect 32845 -8145 32905 -8135
rect 32845 -8185 32855 -8145
rect 32895 -8185 32905 -8145
rect 32845 -8195 32905 -8185
rect 35335 -8145 35395 -8135
rect 35335 -8185 35345 -8145
rect 35385 -8185 35395 -8145
rect 35335 -8195 35395 -8185
rect 37825 -8145 37885 -8135
rect 37825 -8185 37835 -8145
rect 37875 -8185 37885 -8145
rect 37825 -8195 37885 -8185
rect 40315 -8145 40375 -8135
rect 40315 -8185 40325 -8145
rect 40365 -8185 40375 -8145
rect 40315 -8195 40375 -8185
rect 42805 -8145 42865 -8135
rect 42805 -8185 42815 -8145
rect 42855 -8185 42865 -8145
rect 42805 -8195 42865 -8185
rect 45295 -8145 45355 -8135
rect 45295 -8185 45305 -8145
rect 45345 -8185 45355 -8145
rect 45295 -8195 45355 -8185
rect 47785 -8145 47845 -8135
rect 47785 -8185 47795 -8145
rect 47835 -8185 47845 -8145
rect 47785 -8195 47845 -8185
rect 27910 -9345 28190 -9240
rect 7825 -12275 8105 -12185
rect 27910 -12490 28025 -9345
rect 28185 -9640 28255 -9540
rect 7890 -12585 8110 -12495
rect 7890 -12815 7995 -12585
rect 27845 -12595 28190 -12490
rect 7830 -12915 7995 -12815
rect 27855 -12890 28255 -12790
<< via1 >>
rect 1905 6610 1945 6690
rect 30365 -2155 30405 -2145
rect 30365 -2175 30375 -2155
rect 30375 -2175 30395 -2155
rect 30395 -2175 30405 -2155
rect 30365 -2185 30405 -2175
rect 32855 -2155 32895 -2145
rect 32855 -2175 32865 -2155
rect 32865 -2175 32885 -2155
rect 32885 -2175 32895 -2155
rect 32855 -2185 32895 -2175
rect 35345 -2155 35385 -2145
rect 35345 -2175 35355 -2155
rect 35355 -2175 35375 -2155
rect 35375 -2175 35385 -2155
rect 35345 -2185 35385 -2175
rect 37835 -2155 37875 -2145
rect 37835 -2175 37845 -2155
rect 37845 -2175 37865 -2155
rect 37865 -2175 37875 -2155
rect 37835 -2185 37875 -2175
rect 40325 -2155 40365 -2145
rect 40325 -2175 40335 -2155
rect 40335 -2175 40355 -2155
rect 40355 -2175 40365 -2155
rect 40325 -2185 40365 -2175
rect 42815 -2155 42855 -2145
rect 42815 -2175 42825 -2155
rect 42825 -2175 42845 -2155
rect 42845 -2175 42855 -2155
rect 42815 -2185 42855 -2175
rect 45305 -2155 45345 -2145
rect 45305 -2175 45315 -2155
rect 45315 -2175 45335 -2155
rect 45335 -2175 45345 -2155
rect 45305 -2185 45345 -2175
rect 47795 -2155 47835 -2145
rect 47795 -2175 47805 -2155
rect 47805 -2175 47825 -2155
rect 47825 -2175 47835 -2155
rect 47795 -2185 47835 -2175
rect 30365 -8155 30405 -8145
rect 30365 -8175 30375 -8155
rect 30375 -8175 30395 -8155
rect 30395 -8175 30405 -8155
rect 30365 -8185 30405 -8175
rect 32855 -8155 32895 -8145
rect 32855 -8175 32865 -8155
rect 32865 -8175 32885 -8155
rect 32885 -8175 32895 -8155
rect 32855 -8185 32895 -8175
rect 35345 -8155 35385 -8145
rect 35345 -8175 35355 -8155
rect 35355 -8175 35375 -8155
rect 35375 -8175 35385 -8155
rect 35345 -8185 35385 -8175
rect 37835 -8155 37875 -8145
rect 37835 -8175 37845 -8155
rect 37845 -8175 37865 -8155
rect 37865 -8175 37875 -8155
rect 37835 -8185 37875 -8175
rect 40325 -8155 40365 -8145
rect 40325 -8175 40335 -8155
rect 40335 -8175 40355 -8155
rect 40355 -8175 40365 -8155
rect 40325 -8185 40365 -8175
rect 42815 -8155 42855 -8145
rect 42815 -8175 42825 -8155
rect 42825 -8175 42845 -8155
rect 42845 -8175 42855 -8155
rect 42815 -8185 42855 -8175
rect 45305 -8155 45345 -8145
rect 45305 -8175 45315 -8155
rect 45315 -8175 45335 -8155
rect 45335 -8175 45345 -8155
rect 45305 -8185 45345 -8175
rect 47795 -8155 47835 -8145
rect 47795 -8175 47805 -8155
rect 47805 -8175 47825 -8155
rect 47825 -8175 47835 -8155
rect 47795 -8185 47835 -8175
<< metal2 >>
rect 675 6690 4555 6700
rect 675 6610 1905 6690
rect 1945 6610 4555 6690
rect 675 6600 4555 6610
rect 4560 6600 7320 6700
rect 480 -430 615 545
rect 480 -530 4555 -430
rect 4560 -530 7320 -430
rect 28180 -645 28280 600
rect 28185 -1505 28280 -645
rect 30355 -2145 30415 -2135
rect 30355 -2185 30365 -2145
rect 30405 -2185 30415 -2145
rect 480 -7570 615 -6555
rect 480 -7670 4555 -7570
rect 4560 -7670 7320 -7570
rect 30355 -8145 30415 -2185
rect 30355 -8185 30365 -8145
rect 30405 -8185 30415 -8145
rect 30355 -8195 30415 -8185
rect 32845 -2145 32905 -2135
rect 32845 -2185 32855 -2145
rect 32895 -2185 32905 -2145
rect 32845 -8145 32905 -2185
rect 32845 -8185 32855 -8145
rect 32895 -8185 32905 -8145
rect 32845 -8195 32905 -8185
rect 35335 -2145 35395 -2135
rect 35335 -2185 35345 -2145
rect 35385 -2185 35395 -2145
rect 35335 -8145 35395 -2185
rect 35335 -8185 35345 -8145
rect 35385 -8185 35395 -8145
rect 35335 -8195 35395 -8185
rect 37825 -2145 37885 -2135
rect 37825 -2185 37835 -2145
rect 37875 -2185 37885 -2145
rect 37825 -8145 37885 -2185
rect 37825 -8185 37835 -8145
rect 37875 -8185 37885 -8145
rect 37825 -8195 37885 -8185
rect 40315 -2145 40375 -2135
rect 40315 -2185 40325 -2145
rect 40365 -2185 40375 -2145
rect 40315 -8145 40375 -2185
rect 40315 -8185 40325 -8145
rect 40365 -8185 40375 -8145
rect 40315 -8195 40375 -8185
rect 42805 -2145 42865 -2135
rect 42805 -2185 42815 -2145
rect 42855 -2185 42865 -2145
rect 42805 -8145 42865 -2185
rect 42805 -8185 42815 -8145
rect 42855 -8185 42865 -8145
rect 42805 -8195 42865 -8185
rect 45295 -2145 45355 -2135
rect 45295 -2185 45305 -2145
rect 45345 -2185 45355 -2145
rect 45295 -8145 45355 -2185
rect 45295 -8185 45305 -8145
rect 45345 -8185 45355 -8145
rect 45295 -8195 45355 -8185
rect 47785 -2145 47845 -2135
rect 47785 -2185 47795 -2145
rect 47835 -2185 47845 -2145
rect 47785 -8145 47845 -2185
rect 47785 -8185 47795 -8145
rect 47835 -8185 47845 -8145
rect 47785 -8195 47845 -8185
rect 28185 -12275 28285 -10430
use fa_8bit  fa_8bit_0
timestamp 1693914941
transform 1 0 28075 0 1 -3050
box -50 -10 19860 1905
use fa_8bit  fa_8bit_1
timestamp 1693914941
transform 1 0 28075 0 1 -6680
box -50 -10 19860 1905
use fa_8bit  fa_8bit_2
timestamp 1693914941
transform 1 0 8000 0 1 -6685
box -50 -10 19860 1905
use fa_8bit  fa_8bit_3
timestamp 1693914941
transform 1 0 8000 0 1 445
box -50 -10 19860 1905
use fa_8bit  fa_8bit_4
timestamp 1693914941
transform 1 0 28075 0 1 -13820
box -50 -10 19860 1905
use fa_8bit  fa_8bit_5
timestamp 1693914941
transform 1 0 8000 0 1 -13825
box -50 -10 19860 1905
use fa_8bit  fa_8bit_6
timestamp 1693914941
transform 1 0 28075 0 1 450
box -50 -10 19860 1905
use fa_8bit  fa_8bit_7
timestamp 1693914941
transform 1 0 28075 0 1 -10570
box -50 -10 19860 1905
use shifter  shifter_0
timestamp 1693853362
transform 1 0 110 0 1 -740
box -75 -5955 1035 330
use shifter  shifter_1
timestamp 1693853362
transform 1 0 1240 0 1 -740
box -75 -5955 1035 330
use shifter  shifter_2
timestamp 1693853362
transform 1 0 2920 0 1 -740
box -75 -5955 1035 330
use shifter  shifter_3
timestamp 1693853362
transform 1 0 4050 0 1 -740
box -75 -5955 1035 330
use shifter  shifter_4
timestamp 1693853362
transform 1 0 5180 0 1 -740
box -75 -5955 1035 330
use shifter  shifter_5
timestamp 1693853362
transform 1 0 6810 0 1 6390
box -75 -5955 1035 330
use shifter  shifter_6
timestamp 1693853362
transform 1 0 6810 0 1 -740
box -75 -5955 1035 330
use shifter  shifter_7
timestamp 1693853362
transform 1 0 5680 0 1 6390
box -75 -5955 1035 330
use shifter  shifter_8
timestamp 1693853362
transform 1 0 4050 0 1 6390
box -75 -5955 1035 330
use shifter  shifter_9
timestamp 1693853362
transform 1 0 2920 0 1 6390
box -75 -5955 1035 330
use shifter  shifter_10
timestamp 1693853362
transform 1 0 1790 0 1 6390
box -75 -5955 1035 330
use shifter  shifter_11
timestamp 1693853362
transform 1 0 110 0 1 6390
box -75 -5955 1035 330
use shifter  shifter_12
timestamp 1693853362
transform 1 0 6810 0 1 -7880
box -75 -5955 1035 330
use shifter  shifter_13
timestamp 1693853362
transform 1 0 5180 0 1 -7880
box -75 -5955 1035 330
use shifter  shifter_14
timestamp 1693853362
transform 1 0 4050 0 1 -7880
box -75 -5955 1035 330
use shifter  shifter_15
timestamp 1693853362
transform 1 0 2920 0 1 -7880
box -75 -5955 1035 330
use shifter  shifter_16
timestamp 1693853362
transform 1 0 1240 0 1 -7880
box -75 -5955 1035 330
use shifter  shifter_17
timestamp 1693853362
transform 1 0 110 0 1 -7880
box -75 -5955 1035 330
<< end >>
