* NGSPICE file created from and.ext - technology: sky130A

**.subckt and A B VP VN
X0 a_15_n5# B a_15_n300# VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X1 a_225_n300# a_15_n5# VP VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=1.5e+12p ps=9e+06u w=1e+06u l=150000u
X2 a_15_n5# A VP VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_15_n300# A VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1e+12p ps=6e+06u w=1e+06u l=150000u
X4 a_225_n300# a_15_n5# VN VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VP B a_15_n5# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
**.ends


.end
