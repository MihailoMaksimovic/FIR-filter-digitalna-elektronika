magic
tech sky130A
timestamp 1693853362
<< nwell >>
rect 495 310 505 330
rect 485 210 505 310
rect 495 190 505 210
rect 505 -440 1000 -415
rect 90 -555 1000 -440
rect 90 -575 505 -555
rect 485 -1420 1035 -1315
rect 370 -1430 1035 -1420
rect 90 -1455 1035 -1430
rect 90 -1475 505 -1455
rect 495 -2345 740 -2215
rect 90 -2355 740 -2345
rect 90 -2380 505 -2355
rect 500 -3235 735 -3115
rect 90 -3255 735 -3235
rect 90 -3290 505 -3255
rect 500 -4140 720 -4015
rect 90 -4155 720 -4140
rect 90 -4185 505 -4155
rect 495 -5045 735 -4915
rect 90 -5055 735 -5045
rect 90 -5090 505 -5055
<< nmos >>
rect 740 -1730 755 -1630
rect 805 -1730 820 -1630
rect 950 -1730 965 -1630
<< pmos >>
rect 740 -1435 755 -1335
rect 805 -1435 820 -1335
rect 950 -1435 965 -1335
<< ndiff >>
rect 690 -1645 740 -1630
rect 690 -1715 705 -1645
rect 725 -1715 740 -1645
rect 690 -1730 740 -1715
rect 755 -1645 805 -1630
rect 755 -1715 770 -1645
rect 790 -1715 805 -1645
rect 755 -1730 805 -1715
rect 820 -1645 870 -1630
rect 820 -1715 835 -1645
rect 855 -1715 870 -1645
rect 820 -1730 870 -1715
rect 900 -1645 950 -1630
rect 900 -1715 915 -1645
rect 935 -1715 950 -1645
rect 900 -1730 950 -1715
rect 965 -1645 1015 -1630
rect 965 -1715 980 -1645
rect 1000 -1715 1015 -1645
rect 965 -1730 1015 -1715
<< pdiff >>
rect 690 -1350 740 -1335
rect 690 -1420 705 -1350
rect 725 -1420 740 -1350
rect 690 -1435 740 -1420
rect 755 -1350 805 -1335
rect 755 -1420 770 -1350
rect 790 -1420 805 -1350
rect 755 -1435 805 -1420
rect 820 -1350 870 -1335
rect 820 -1420 835 -1350
rect 855 -1420 870 -1350
rect 820 -1435 870 -1420
rect 900 -1350 950 -1335
rect 900 -1420 915 -1350
rect 935 -1420 950 -1350
rect 900 -1435 950 -1420
rect 965 -1350 1015 -1335
rect 965 -1420 980 -1350
rect 1000 -1420 1015 -1350
rect 965 -1435 1015 -1420
<< ndiffc >>
rect 705 -1715 725 -1645
rect 770 -1715 790 -1645
rect 835 -1715 855 -1645
rect 915 -1715 935 -1645
rect 980 -1715 1000 -1645
<< pdiffc >>
rect 705 -1420 725 -1350
rect 770 -1420 790 -1350
rect 835 -1420 855 -1350
rect 915 -1420 935 -1350
rect 980 -1420 1000 -1350
<< psubdiff >>
rect 640 -1645 690 -1630
rect 640 -1715 655 -1645
rect 675 -1715 690 -1645
rect 640 -1730 690 -1715
<< nsubdiff >>
rect 640 -1350 690 -1335
rect 640 -1420 655 -1350
rect 675 -1420 690 -1350
rect 640 -1435 690 -1420
<< psubdiffcont >>
rect 655 -1715 675 -1645
<< nsubdiffcont >>
rect 655 -1420 675 -1350
<< poly >>
rect -75 180 -35 190
rect -75 160 -65 180
rect -45 160 -35 180
rect -75 150 -35 160
rect -50 -810 -35 150
rect -10 -310 30 -300
rect -10 -330 0 -310
rect 20 -330 30 -310
rect -10 -340 30 -330
rect -75 -820 -35 -810
rect -75 -840 -65 -820
rect -45 -840 -35 -820
rect -75 -850 -35 -840
rect -50 -1730 -35 -850
rect 15 -1200 30 -340
rect 480 -385 520 -375
rect 480 -405 490 -385
rect 510 -400 520 -385
rect 590 -385 630 -375
rect 590 -400 600 -385
rect 510 -405 600 -400
rect 620 -405 630 -385
rect 480 -415 630 -405
rect 90 -720 130 -710
rect 90 -740 100 -720
rect 120 -740 130 -720
rect 90 -750 130 -740
rect 480 -720 605 -710
rect 480 -740 490 -720
rect 510 -725 605 -720
rect 510 -740 520 -725
rect 480 -750 520 -740
rect 90 -830 105 -750
rect 90 -840 130 -830
rect 90 -860 100 -840
rect 120 -860 130 -840
rect 90 -870 130 -860
rect -10 -1210 30 -1200
rect -10 -1230 0 -1210
rect 20 -1230 30 -1210
rect -10 -1240 30 -1230
rect -75 -1740 -35 -1730
rect -75 -1760 -65 -1740
rect -45 -1760 -35 -1740
rect -75 -1770 -35 -1760
rect -50 -2630 -35 -1770
rect 15 -2100 30 -1240
rect 590 -1275 605 -725
rect 590 -1285 630 -1275
rect 590 -1305 600 -1285
rect 620 -1305 630 -1285
rect 590 -1315 630 -1305
rect 740 -1335 755 -1320
rect 805 -1335 820 -1320
rect 950 -1335 965 -1320
rect 740 -1455 755 -1435
rect 715 -1465 755 -1455
rect 715 -1485 725 -1465
rect 745 -1485 755 -1465
rect 715 -1495 755 -1485
rect 90 -1620 130 -1610
rect 90 -1640 100 -1620
rect 120 -1640 130 -1620
rect 90 -1650 130 -1640
rect 480 -1620 605 -1610
rect 480 -1640 490 -1620
rect 510 -1625 605 -1620
rect 510 -1640 520 -1625
rect 480 -1650 520 -1640
rect 90 -1730 105 -1650
rect 90 -1740 130 -1730
rect 90 -1760 100 -1740
rect 120 -1760 130 -1740
rect 90 -1770 130 -1760
rect -10 -2110 30 -2100
rect -10 -2130 0 -2110
rect 20 -2130 30 -2110
rect -10 -2140 30 -2130
rect -75 -2640 -35 -2630
rect -75 -2660 -65 -2640
rect -45 -2660 -35 -2640
rect -75 -2670 -35 -2660
rect -50 -3530 -35 -2670
rect 15 -3000 30 -2140
rect 590 -2175 605 -1625
rect 740 -1630 755 -1495
rect 805 -1530 820 -1435
rect 950 -1455 965 -1435
rect 925 -1465 965 -1455
rect 925 -1485 935 -1465
rect 955 -1485 965 -1465
rect 925 -1495 965 -1485
rect 780 -1540 820 -1530
rect 780 -1560 790 -1540
rect 810 -1560 820 -1540
rect 780 -1570 820 -1560
rect 805 -1630 820 -1570
rect 950 -1630 965 -1495
rect 740 -1745 755 -1730
rect 805 -1745 820 -1730
rect 950 -1745 965 -1730
rect 590 -2185 630 -2175
rect 590 -2205 600 -2185
rect 620 -2205 630 -2185
rect 590 -2215 630 -2205
rect 90 -2520 130 -2510
rect 90 -2540 100 -2520
rect 120 -2540 130 -2520
rect 90 -2550 130 -2540
rect 460 -2520 605 -2510
rect 460 -2540 470 -2520
rect 490 -2525 605 -2520
rect 490 -2540 500 -2525
rect 460 -2550 500 -2540
rect 90 -2630 105 -2550
rect 90 -2640 130 -2630
rect 90 -2660 100 -2640
rect 120 -2660 130 -2640
rect 90 -2670 130 -2660
rect -10 -3010 30 -3000
rect -10 -3030 0 -3010
rect 20 -3030 30 -3010
rect -10 -3040 30 -3030
rect -75 -3540 -35 -3530
rect -75 -3560 -65 -3540
rect -45 -3560 -35 -3540
rect -75 -3570 -35 -3560
rect -50 -4430 -35 -3570
rect -75 -4440 -35 -4430
rect -75 -4460 -65 -4440
rect -45 -4460 -35 -4440
rect -75 -4470 -35 -4460
rect -50 -5330 -35 -4470
rect -75 -5340 -35 -5330
rect -75 -5360 -65 -5340
rect -45 -5360 -35 -5340
rect -75 -5370 -35 -5360
rect 15 -3900 30 -3040
rect 590 -3075 605 -2525
rect 590 -3085 630 -3075
rect 590 -3105 600 -3085
rect 620 -3105 630 -3085
rect 590 -3115 630 -3105
rect 90 -3420 130 -3410
rect 90 -3440 100 -3420
rect 120 -3440 130 -3420
rect 90 -3450 130 -3440
rect 460 -3420 605 -3410
rect 460 -3440 470 -3420
rect 490 -3425 605 -3420
rect 490 -3440 500 -3425
rect 460 -3450 500 -3440
rect 90 -3530 105 -3450
rect 90 -3540 130 -3530
rect 90 -3560 100 -3540
rect 120 -3560 130 -3540
rect 90 -3570 130 -3560
rect 15 -3910 55 -3900
rect 15 -3930 25 -3910
rect 45 -3930 55 -3910
rect 15 -3940 55 -3930
rect 15 -4800 30 -3940
rect 590 -3975 605 -3425
rect 590 -3985 630 -3975
rect 590 -4005 600 -3985
rect 620 -4005 630 -3985
rect 590 -4015 630 -4005
rect 90 -4320 130 -4310
rect 90 -4340 100 -4320
rect 120 -4340 130 -4320
rect 90 -4350 130 -4340
rect 460 -4320 605 -4310
rect 460 -4340 470 -4320
rect 490 -4325 605 -4320
rect 490 -4340 500 -4325
rect 460 -4350 500 -4340
rect 90 -4430 105 -4350
rect 90 -4440 130 -4430
rect 90 -4460 100 -4440
rect 120 -4460 130 -4440
rect 90 -4470 130 -4460
rect 15 -4810 55 -4800
rect 15 -4830 25 -4810
rect 45 -4830 55 -4810
rect 15 -4840 55 -4830
rect 15 -5700 30 -4840
rect 590 -4875 605 -4325
rect 590 -4885 630 -4875
rect 590 -4905 600 -4885
rect 620 -4905 630 -4885
rect 590 -4915 630 -4905
rect 90 -5220 130 -5210
rect 90 -5240 100 -5220
rect 120 -5240 130 -5220
rect 90 -5250 130 -5240
rect 460 -5220 605 -5210
rect 460 -5240 470 -5220
rect 490 -5225 605 -5220
rect 490 -5240 500 -5225
rect 460 -5250 500 -5240
rect 90 -5330 105 -5250
rect 90 -5340 130 -5330
rect 90 -5360 100 -5340
rect 120 -5360 130 -5340
rect 90 -5370 130 -5360
rect 590 -5345 605 -5225
rect 590 -5355 630 -5345
rect 590 -5375 600 -5355
rect 620 -5375 630 -5355
rect 590 -5385 630 -5375
rect 15 -5710 55 -5700
rect 15 -5730 25 -5710
rect 45 -5730 55 -5710
rect 15 -5740 55 -5730
<< polycont >>
rect -65 160 -45 180
rect 0 -330 20 -310
rect -65 -840 -45 -820
rect 490 -405 510 -385
rect 600 -405 620 -385
rect 100 -740 120 -720
rect 490 -740 510 -720
rect 100 -860 120 -840
rect 0 -1230 20 -1210
rect -65 -1760 -45 -1740
rect 600 -1305 620 -1285
rect 725 -1485 745 -1465
rect 100 -1640 120 -1620
rect 490 -1640 510 -1620
rect 100 -1760 120 -1740
rect 0 -2130 20 -2110
rect -65 -2660 -45 -2640
rect 935 -1485 955 -1465
rect 790 -1560 810 -1540
rect 600 -2205 620 -2185
rect 100 -2540 120 -2520
rect 470 -2540 490 -2520
rect 100 -2660 120 -2640
rect 0 -3030 20 -3010
rect -65 -3560 -45 -3540
rect -65 -4460 -45 -4440
rect -65 -5360 -45 -5340
rect 600 -3105 620 -3085
rect 100 -3440 120 -3420
rect 470 -3440 490 -3420
rect 100 -3560 120 -3540
rect 25 -3930 45 -3910
rect 600 -4005 620 -3985
rect 100 -4340 120 -4320
rect 470 -4340 490 -4320
rect 100 -4460 120 -4440
rect 25 -4830 45 -4810
rect 600 -4905 620 -4885
rect 100 -5240 120 -5220
rect 470 -5240 490 -5220
rect 100 -5360 120 -5340
rect 600 -5375 620 -5355
rect 25 -5730 45 -5710
<< locali >>
rect -75 180 100 190
rect -75 160 -65 180
rect -45 170 100 180
rect 495 170 570 190
rect -45 160 -35 170
rect -75 150 -35 160
rect -10 -310 30 -300
rect -10 -330 0 -310
rect 20 -320 30 -310
rect 20 -330 110 -320
rect -10 -340 110 -330
rect 480 -385 520 -375
rect 35 -415 125 -395
rect 480 -405 490 -385
rect 510 -405 520 -385
rect 480 -415 520 -405
rect 35 -785 55 -415
rect 550 -555 570 170
rect 590 -385 630 -375
rect 590 -405 600 -385
rect 620 -395 630 -385
rect 620 -405 1035 -395
rect 590 -415 1035 -405
rect 550 -575 640 -555
rect 550 -650 625 -630
rect 630 -645 645 -630
rect 90 -720 130 -710
rect 90 -740 100 -720
rect 120 -740 130 -720
rect 90 -750 130 -740
rect 460 -720 520 -710
rect 460 -740 490 -720
rect 510 -740 520 -720
rect 460 -750 520 -740
rect 35 -805 125 -785
rect -75 -820 -35 -810
rect -75 -840 -65 -820
rect -45 -830 -35 -820
rect -45 -840 130 -830
rect -75 -850 100 -840
rect 90 -860 100 -850
rect 120 -860 130 -840
rect 90 -870 130 -860
rect -10 -1210 30 -1200
rect -10 -1230 0 -1210
rect 20 -1220 30 -1210
rect 20 -1230 115 -1220
rect -10 -1240 115 -1230
rect 550 -1295 570 -650
rect 35 -1315 110 -1295
rect 505 -1315 570 -1295
rect 590 -1285 630 -1275
rect 590 -1305 600 -1285
rect 620 -1305 630 -1285
rect 590 -1315 630 -1305
rect 35 -1685 55 -1315
rect 590 -1455 610 -1315
rect 645 -1350 735 -1340
rect 645 -1420 655 -1350
rect 675 -1420 705 -1350
rect 725 -1420 735 -1350
rect 645 -1430 735 -1420
rect 760 -1350 800 -1340
rect 760 -1420 770 -1350
rect 790 -1420 800 -1350
rect 760 -1430 800 -1420
rect 825 -1350 865 -1340
rect 825 -1420 835 -1350
rect 855 -1420 865 -1350
rect 825 -1430 865 -1420
rect 905 -1350 945 -1340
rect 905 -1420 915 -1350
rect 935 -1420 945 -1350
rect 905 -1430 945 -1420
rect 970 -1350 1010 -1340
rect 970 -1420 980 -1350
rect 1000 -1420 1010 -1350
rect 970 -1430 1010 -1420
rect 845 -1455 865 -1430
rect 990 -1455 1010 -1430
rect 590 -1465 755 -1455
rect 590 -1475 725 -1465
rect 715 -1485 725 -1475
rect 745 -1485 755 -1465
rect 715 -1495 755 -1485
rect 845 -1465 965 -1455
rect 845 -1475 935 -1465
rect 545 -1540 820 -1530
rect 545 -1550 790 -1540
rect 90 -1620 130 -1610
rect 90 -1640 100 -1620
rect 120 -1640 130 -1620
rect 90 -1650 130 -1640
rect 480 -1620 520 -1610
rect 480 -1640 490 -1620
rect 510 -1640 520 -1620
rect 480 -1650 520 -1640
rect 35 -1705 100 -1685
rect -75 -1740 -35 -1730
rect -75 -1760 -65 -1740
rect -45 -1750 -35 -1740
rect 90 -1740 130 -1730
rect 90 -1750 100 -1740
rect -45 -1760 100 -1750
rect 120 -1760 130 -1740
rect -75 -1770 130 -1760
rect -10 -2110 30 -2100
rect -10 -2130 0 -2110
rect 20 -2120 30 -2110
rect 20 -2130 160 -2120
rect -10 -2140 160 -2130
rect 545 -2195 565 -1550
rect 780 -1560 790 -1550
rect 810 -1560 820 -1540
rect 780 -1570 820 -1560
rect 845 -1595 865 -1475
rect 925 -1485 935 -1475
rect 955 -1485 965 -1465
rect 925 -1495 965 -1485
rect 990 -1475 1035 -1455
rect 780 -1615 865 -1595
rect 780 -1635 800 -1615
rect 925 -1635 945 -1630
rect 990 -1635 1010 -1475
rect 645 -1645 735 -1635
rect 645 -1715 655 -1645
rect 675 -1715 705 -1645
rect 725 -1715 735 -1645
rect 645 -1725 735 -1715
rect 760 -1645 800 -1635
rect 760 -1715 770 -1645
rect 790 -1715 800 -1645
rect 760 -1725 800 -1715
rect 825 -1645 865 -1635
rect 825 -1715 835 -1645
rect 855 -1715 865 -1645
rect 825 -1725 865 -1715
rect 905 -1645 945 -1635
rect 905 -1715 915 -1645
rect 935 -1715 945 -1645
rect 905 -1725 945 -1715
rect 970 -1645 1010 -1635
rect 970 -1715 980 -1645
rect 1000 -1715 1010 -1645
rect 970 -1725 1010 -1715
rect 35 -2215 120 -2195
rect 505 -2215 565 -2195
rect 590 -2185 630 -2175
rect 590 -2205 600 -2185
rect 620 -2205 630 -2185
rect 590 -2215 630 -2205
rect 35 -2585 55 -2215
rect 590 -2355 610 -2215
rect 590 -2375 635 -2355
rect 545 -2450 645 -2430
rect 90 -2520 130 -2510
rect 90 -2540 100 -2520
rect 120 -2540 130 -2520
rect 90 -2550 130 -2540
rect 460 -2520 500 -2510
rect 460 -2540 470 -2520
rect 490 -2540 500 -2520
rect 460 -2550 500 -2540
rect 35 -2605 120 -2585
rect -75 -2640 -35 -2630
rect -75 -2660 -65 -2640
rect -45 -2650 -35 -2640
rect 90 -2640 130 -2630
rect 90 -2650 100 -2640
rect -45 -2660 100 -2650
rect 120 -2660 130 -2640
rect -75 -2670 130 -2660
rect -10 -3010 30 -3000
rect -10 -3030 0 -3010
rect 20 -3020 30 -3010
rect 20 -3030 180 -3020
rect -10 -3040 180 -3030
rect 545 -3095 565 -2450
rect 35 -3115 115 -3095
rect 505 -3115 565 -3095
rect 590 -3085 630 -3075
rect 590 -3105 600 -3085
rect 620 -3105 630 -3085
rect 590 -3115 630 -3105
rect 35 -3485 55 -3115
rect 590 -3255 610 -3115
rect 590 -3275 630 -3255
rect 545 -3350 625 -3330
rect 90 -3420 130 -3410
rect 90 -3440 100 -3420
rect 120 -3440 130 -3420
rect 90 -3450 130 -3440
rect 460 -3420 500 -3410
rect 460 -3440 470 -3420
rect 490 -3440 500 -3420
rect 460 -3450 500 -3440
rect 35 -3505 110 -3485
rect -75 -3540 -35 -3530
rect -75 -3560 -65 -3540
rect -45 -3550 -35 -3540
rect 90 -3540 130 -3530
rect 90 -3550 100 -3540
rect -45 -3560 100 -3550
rect 120 -3560 130 -3540
rect -75 -3570 130 -3560
rect 15 -3910 55 -3900
rect 15 -3930 25 -3910
rect 45 -3920 55 -3910
rect 45 -3930 170 -3920
rect 15 -3940 170 -3930
rect 545 -3995 565 -3350
rect 35 -4015 120 -3995
rect 500 -4015 565 -3995
rect 590 -3985 630 -3975
rect 590 -4005 600 -3985
rect 620 -4005 630 -3985
rect 590 -4015 630 -4005
rect 35 -4385 55 -4015
rect 590 -4155 610 -4015
rect 590 -4175 630 -4155
rect 545 -4250 625 -4230
rect 90 -4320 130 -4310
rect 90 -4340 100 -4320
rect 120 -4340 130 -4320
rect 90 -4350 130 -4340
rect 460 -4320 500 -4310
rect 460 -4340 470 -4320
rect 490 -4340 500 -4320
rect 460 -4350 500 -4340
rect 35 -4405 115 -4385
rect -75 -4440 -35 -4430
rect -75 -4460 -65 -4440
rect -45 -4450 -35 -4440
rect 90 -4440 130 -4430
rect 90 -4450 100 -4440
rect -45 -4460 100 -4450
rect 120 -4460 130 -4440
rect -75 -4470 130 -4460
rect 15 -4810 55 -4800
rect 15 -4830 25 -4810
rect 45 -4820 55 -4810
rect 45 -4830 175 -4820
rect 15 -4840 175 -4830
rect 545 -4895 565 -4250
rect 35 -4915 115 -4895
rect 505 -4915 565 -4895
rect 590 -4885 630 -4875
rect 590 -4905 600 -4885
rect 620 -4905 630 -4885
rect 590 -4915 630 -4905
rect 35 -5285 55 -4915
rect 590 -5055 610 -4915
rect 590 -5075 635 -5055
rect 545 -5150 635 -5130
rect 90 -5220 130 -5210
rect 90 -5240 100 -5220
rect 120 -5240 130 -5220
rect 90 -5250 130 -5240
rect 460 -5220 500 -5210
rect 460 -5240 470 -5220
rect 490 -5240 500 -5220
rect 460 -5250 500 -5240
rect 35 -5305 110 -5285
rect -75 -5340 -35 -5330
rect -75 -5360 -65 -5340
rect -45 -5350 -35 -5340
rect 90 -5340 130 -5330
rect 90 -5350 100 -5340
rect -45 -5360 100 -5350
rect 120 -5360 130 -5340
rect -75 -5370 130 -5360
rect 15 -5710 55 -5700
rect 15 -5730 25 -5710
rect 45 -5720 55 -5710
rect 45 -5730 170 -5720
rect 15 -5740 170 -5730
rect 545 -5795 565 -5150
rect 590 -5355 630 -5345
rect 590 -5375 600 -5355
rect 620 -5365 630 -5355
rect 620 -5375 1035 -5365
rect 590 -5385 1035 -5375
rect 495 -5815 565 -5795
<< viali >>
rect 655 -1420 675 -1350
rect 705 -1420 725 -1350
rect 915 -1420 935 -1350
rect 655 -1715 675 -1645
rect 705 -1715 725 -1645
rect 835 -1715 855 -1645
rect 915 -1715 935 -1645
<< metal1 >>
rect 500 -65 570 15
rect 495 -235 570 -65
rect 505 -240 570 -235
rect 535 -730 570 -240
rect 535 -780 620 -730
rect 535 -885 570 -780
rect 500 -980 570 -885
rect 505 -985 570 -980
rect 535 -1040 570 -985
rect 500 -1130 570 -1040
rect 505 -1140 570 -1130
rect 535 -1630 570 -1140
rect 620 -1345 1030 -1335
rect 620 -1425 645 -1345
rect 685 -1350 1030 -1345
rect 685 -1420 705 -1350
rect 725 -1420 915 -1350
rect 935 -1420 1030 -1350
rect 685 -1425 1030 -1420
rect 620 -1435 1030 -1425
rect 535 -1645 1030 -1630
rect 535 -1680 655 -1645
rect 535 -1785 570 -1680
rect 620 -1715 655 -1680
rect 675 -1715 705 -1645
rect 725 -1715 835 -1645
rect 855 -1715 915 -1645
rect 935 -1715 1030 -1645
rect 620 -1730 1030 -1715
rect 505 -1885 570 -1785
rect 535 -1940 570 -1885
rect 495 -2040 570 -1940
rect 535 -2530 570 -2040
rect 535 -2630 635 -2530
rect 535 -2685 570 -2630
rect 495 -2785 570 -2685
rect 535 -2840 570 -2785
rect 490 -2940 570 -2840
rect 535 -3430 570 -2940
rect 535 -3530 635 -3430
rect 535 -3585 570 -3530
rect 495 -3685 570 -3585
rect 535 -3740 570 -3685
rect 495 -3840 570 -3740
rect 535 -4330 570 -3840
rect 535 -4430 635 -4330
rect 535 -4485 570 -4430
rect 490 -4585 570 -4485
rect 535 -4640 570 -4585
rect 495 -4740 570 -4640
rect 535 -5230 570 -4740
rect 535 -5330 635 -5230
rect 535 -5385 570 -5330
rect 495 -5485 570 -5385
rect 535 -5540 570 -5485
rect 490 -5640 570 -5540
<< via1 >>
rect 380 225 415 295
rect 375 -525 420 -445
rect 375 -680 415 -600
rect 645 -525 685 -445
rect 375 -1420 420 -1340
rect 375 -1575 415 -1495
rect 645 -1350 685 -1345
rect 645 -1420 655 -1350
rect 655 -1420 675 -1350
rect 675 -1420 685 -1350
rect 645 -1425 685 -1420
rect 375 -2325 415 -2245
rect 375 -2480 415 -2400
rect 645 -2325 685 -2245
rect 375 -3225 415 -3145
rect 375 -3380 415 -3300
rect 645 -3225 685 -3145
rect 375 -4125 415 -4045
rect 375 -4280 415 -4200
rect 645 -4125 685 -4045
rect 375 -5025 415 -4945
rect 375 -5180 415 -5100
rect 645 -5025 685 -4945
rect 375 -5925 415 -5845
<< metal2 >>
rect 370 295 570 310
rect 370 225 380 295
rect 415 225 570 295
rect 370 210 570 225
rect 530 -435 570 210
rect 370 -445 690 -435
rect 370 -525 375 -445
rect 420 -525 645 -445
rect 685 -525 690 -445
rect 370 -535 690 -525
rect 530 -590 570 -535
rect 370 -600 570 -590
rect 370 -680 375 -600
rect 415 -680 570 -600
rect 370 -690 570 -680
rect 530 -1335 570 -690
rect 370 -1340 690 -1335
rect 370 -1420 375 -1340
rect 420 -1345 690 -1340
rect 420 -1420 645 -1345
rect 370 -1425 645 -1420
rect 685 -1425 690 -1345
rect 370 -1435 690 -1425
rect 530 -1490 570 -1435
rect 370 -1495 570 -1490
rect 370 -1575 375 -1495
rect 415 -1575 570 -1495
rect 370 -1590 570 -1575
rect 530 -2235 570 -1590
rect 370 -2245 740 -2235
rect 370 -2325 375 -2245
rect 415 -2325 645 -2245
rect 685 -2325 740 -2245
rect 370 -2335 740 -2325
rect 530 -2390 570 -2335
rect 370 -2400 570 -2390
rect 370 -2480 375 -2400
rect 415 -2480 570 -2400
rect 370 -2490 570 -2480
rect 530 -3135 570 -2490
rect 370 -3145 740 -3135
rect 370 -3225 375 -3145
rect 415 -3225 645 -3145
rect 685 -3225 740 -3145
rect 370 -3235 740 -3225
rect 530 -3290 570 -3235
rect 370 -3300 570 -3290
rect 370 -3380 375 -3300
rect 415 -3380 570 -3300
rect 370 -3390 570 -3380
rect 530 -4035 570 -3390
rect 370 -4045 740 -4035
rect 370 -4125 375 -4045
rect 415 -4125 645 -4045
rect 685 -4125 740 -4045
rect 370 -4135 740 -4125
rect 530 -4190 570 -4135
rect 370 -4200 570 -4190
rect 370 -4280 375 -4200
rect 415 -4280 570 -4200
rect 370 -4290 570 -4280
rect 530 -4935 570 -4290
rect 370 -4945 740 -4935
rect 370 -5025 375 -4945
rect 415 -5025 645 -4945
rect 685 -5025 740 -4945
rect 370 -5035 740 -5025
rect 530 -5090 570 -5035
rect 370 -5100 570 -5090
rect 370 -5180 375 -5100
rect 415 -5180 570 -5100
rect 370 -5190 570 -5180
rect 530 -5835 570 -5190
rect 370 -5845 570 -5835
rect 370 -5925 375 -5845
rect 415 -5925 570 -5845
rect 370 -5935 570 -5925
use and  and_0
timestamp 1693223098
transform 1 0 210 0 1 215
box -120 -315 295 115
use and  and_1
timestamp 1693223098
transform 1 0 210 0 -1 -440
box -120 -315 295 115
use and  and_2
timestamp 1693223098
transform 1 0 210 0 1 -685
box -120 -315 295 115
use and  and_3
timestamp 1693223098
transform 1 0 210 0 -1 -1340
box -120 -315 295 115
use and  and_4
timestamp 1693223098
transform 1 0 210 0 1 -1585
box -120 -315 295 115
use and  and_5
timestamp 1693223098
transform 1 0 210 0 -1 -2240
box -120 -315 295 115
use and  and_6
timestamp 1693223098
transform 1 0 210 0 1 -2485
box -120 -315 295 115
use and  and_7
timestamp 1693223098
transform 1 0 210 0 -1 -3140
box -120 -315 295 115
use and  and_8
timestamp 1693223098
transform 1 0 210 0 1 -3385
box -120 -315 295 115
use and  and_9
timestamp 1693223098
transform 1 0 210 0 -1 -4040
box -120 -315 295 115
use and  and_10
timestamp 1693223098
transform 1 0 210 0 1 -4285
box -120 -315 295 115
use and  and_11
timestamp 1693223098
transform 1 0 210 0 -1 -4940
box -120 -315 295 115
use and  and_12
timestamp 1693223098
transform 1 0 210 0 1 -5185
box -120 -315 295 115
use and  and_13
timestamp 1693223098
transform 1 0 210 0 -1 -5840
box -120 -315 295 115
use or  or_0
timestamp 1693223168
transform 1 0 740 0 1 -530
box -120 -315 295 115
use or  or_1
timestamp 1693223168
transform 1 0 740 0 1 -2330
box -120 -315 295 115
use or  or_2
timestamp 1693223168
transform 1 0 740 0 1 -3230
box -120 -315 295 115
use or  or_3
timestamp 1693223168
transform 1 0 740 0 1 -4130
box -120 -315 295 115
use or  or_4
timestamp 1693223168
transform 1 0 740 0 1 -5030
box -120 -315 295 115
<< labels >>
rlabel metal1 620 -1680 620 -1680 7 VN
port 5 w
rlabel metal1 620 -1385 620 -1385 7 VP
port 4 w
rlabel locali 1035 -1465 1035 -1465 3 X
port 3 e
<< end >>
