magic
tech sky130A
timestamp 1693913107
<< nwell >>
rect 1110 290 1215 430
rect 0 -420 275 -385
rect 0 -505 415 -420
<< poly >>
rect -15 800 25 810
rect -15 780 -5 800
rect 15 780 25 800
rect -15 770 25 780
rect -95 760 -55 770
rect -95 740 -85 760
rect -65 740 -55 760
rect -95 730 -55 740
rect -15 -200 0 770
rect 850 -50 890 -40
rect 850 -70 860 -50
rect 880 -70 890 -50
rect 850 -80 890 -70
rect -15 -210 25 -200
rect -15 -230 -5 -210
rect 15 -230 25 -210
rect -15 -240 25 -230
rect 410 -210 450 -200
rect 410 -230 420 -210
rect 440 -230 450 -210
rect 410 -240 450 -230
rect -15 -285 25 -275
rect -15 -305 -5 -285
rect 15 -305 25 -285
rect -15 -315 25 -305
rect -80 -605 -40 -595
rect -80 -625 -70 -605
rect -50 -625 -40 -605
rect -80 -635 -40 -625
rect -15 -890 0 -315
rect 410 -595 425 -240
rect 850 -435 865 -80
rect 850 -445 890 -435
rect 850 -465 860 -445
rect 880 -465 890 -445
rect 850 -475 890 -465
rect 410 -605 450 -595
rect 410 -625 420 -605
rect 440 -625 450 -605
rect 410 -635 450 -625
rect -40 -900 0 -890
rect -40 -920 -30 -900
rect -10 -920 0 -900
rect -40 -930 0 -920
<< polycont >>
rect -5 780 15 800
rect -85 740 -65 760
rect 860 -70 880 -50
rect -5 -230 15 -210
rect 420 -230 440 -210
rect -5 -305 15 -285
rect -70 -625 -50 -605
rect 860 -465 880 -445
rect 420 -625 440 -605
rect -30 -920 -10 -900
<< locali >>
rect -15 955 985 975
rect -15 810 5 955
rect -15 800 25 810
rect -15 780 -5 800
rect 15 780 25 800
rect -15 770 25 780
rect -95 760 -55 770
rect -95 740 -85 760
rect -65 750 -55 760
rect 965 750 985 955
rect -65 740 0 750
rect -95 730 0 740
rect 965 730 1215 750
rect -95 -440 -75 730
rect 1160 280 1175 290
rect 1155 135 1175 280
rect -140 -460 -75 -440
rect -55 115 0 135
rect 1155 115 1190 135
rect -140 -690 -120 -460
rect -55 -480 -35 115
rect 1155 -40 1175 115
rect 850 -50 1175 -40
rect 850 -70 860 -50
rect 880 -60 1175 -50
rect 880 -70 890 -60
rect 850 -80 890 -70
rect -15 -210 25 -200
rect -15 -230 -5 -210
rect 15 -230 25 -210
rect -15 -240 25 -230
rect 410 -210 450 -200
rect 410 -230 420 -210
rect 440 -230 450 -210
rect 410 -240 450 -230
rect -15 -285 25 -275
rect -15 -305 -5 -285
rect 15 -305 25 -285
rect -15 -315 25 -305
rect 820 -315 890 -295
rect 850 -445 890 -435
rect 850 -455 860 -445
rect -60 -500 -35 -480
rect 470 -465 860 -455
rect 880 -465 890 -445
rect 470 -475 890 -465
rect -60 -595 -40 -500
rect -80 -605 -40 -595
rect -80 -625 -70 -605
rect -50 -615 -40 -605
rect 410 -605 450 -595
rect -50 -625 20 -615
rect -80 -635 20 -625
rect 410 -625 420 -605
rect 440 -625 450 -605
rect 410 -635 450 -625
rect -140 -710 25 -690
rect -40 -900 0 -890
rect -40 -920 -30 -900
rect -10 -910 0 -900
rect 470 -910 490 -475
rect -10 -920 490 -910
rect -40 -930 490 -920
<< metal1 >>
rect 1140 20 1255 115
rect 70 -45 685 20
rect 1155 15 1255 20
<< via1 >>
rect 770 320 810 400
rect 75 160 115 240
rect 25 -130 65 -50
rect 75 -130 115 -50
rect 700 -425 740 -345
rect 25 -880 65 -800
<< metal2 >>
rect 695 400 825 410
rect 695 320 770 400
rect 810 320 825 400
rect 20 240 120 250
rect 20 160 75 240
rect 115 160 120 240
rect 20 -50 120 160
rect 20 -130 25 -50
rect 65 -130 75 -50
rect 115 -130 120 -50
rect 20 -800 120 -130
rect 695 -345 825 320
rect 695 -425 700 -345
rect 740 -425 825 -345
rect 695 -435 825 -425
rect 20 -880 25 -800
rect 65 -880 120 -800
rect 20 -890 120 -880
use and  and_0
timestamp 1693223098
transform 1 0 120 0 -1 -340
box -120 -315 295 115
use and  and_1
timestamp 1693223098
transform 1 0 120 0 1 -590
box -120 -315 295 115
use or  or_0
timestamp 1693223168
transform 1 0 535 0 -1 -340
box -120 -315 295 115
use xor_  xor__0
timestamp 1693670599
transform 1 0 275 0 1 0
box -275 0 885 875
use xor_  xor__1
timestamp 1693670599
transform 1 0 1455 0 1 0
box -275 0 885 875
<< end >>
